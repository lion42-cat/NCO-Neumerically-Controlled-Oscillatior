`timescale 1ns / 1fs
//////////////////////////////////////////////////////////////////////////////////
module sin_cos_rom(clk, rst, addr_in, sin_out, cos_out);
input clk,rst;
input [15:0] addr_in;
output [15:0] sin_out, cos_out;

wire [15:0] addr;
reg [14:0] addr_rom; //{1'b0, addr[13:0]} //주소 음수 표현 방지
reg [31:0] data_rom;
reg [15:0] sin_out, cos_out;
//in
	dff_16bit rom_a(addr_in, clk, rst, addr);

//calculate
	//n사분면 bit에 따라 address_rom 조절
	always @ (addr)
		begin
			case(addr[15:14])
				2'b00 : addr_rom <= {1'b0, addr[13:0]};
				2'b01 : addr_rom <= {1'b0, (14'd16383 - addr[13:0])}; //맨 앞자리인 14번째 bit는 부호 bit임. 
							     						          //2^14-1 - addr[13:0]
				2'b10 : addr_rom <= {1'b0, addr[13:0]};
				2'b11 : addr_rom <= {1'b0, (14'd16383 - addr[13:0])};
				default : addr_rom <= 2'b11000011110000;
			endcase
		end
		
	always @ (addr_rom) //addr_rom은 13bit임!! (n사분면 bit 없음)
		begin
			case (addr_rom)
                15'd0 : data_rom <= {16'd0, 16'd32767};
                15'd1 : data_rom <= {16'd3, 16'd32767};
                15'd2 : data_rom <= {16'd6, 16'd32767};
                15'd3 : data_rom <= {16'd9, 16'd32767};
                15'd4 : data_rom <= {16'd12, 16'd32767};
                15'd5 : data_rom <= {16'd15, 16'd32767};
                15'd6 : data_rom <= {16'd18, 16'd32767};
                15'd7 : data_rom <= {16'd21, 16'd32767};
                15'd8 : data_rom <= {16'd25, 16'd32767};
                15'd9 : data_rom <= {16'd28, 16'd32767};
                15'd10 : data_rom <= {16'd31, 16'd32767};
                15'd11 : data_rom <= {16'd34, 16'd32767};
                15'd12 : data_rom <= {16'd37, 16'd32767};
                15'd13 : data_rom <= {16'd40, 16'd32767};
                15'd14 : data_rom <= {16'd43, 16'd32767};
                15'd15 : data_rom <= {16'd47, 16'd32767};
                15'd16 : data_rom <= {16'd50, 16'd32767};
                15'd17 : data_rom <= {16'd53, 16'd32767};
                15'd18 : data_rom <= {16'd56, 16'd32767};
                15'd19 : data_rom <= {16'd59, 16'd32767};
                15'd20 : data_rom <= {16'd62, 16'd32767};
                15'd21 : data_rom <= {16'd65, 16'd32767};
                15'd22 : data_rom <= {16'd69, 16'd32767};
                15'd23 : data_rom <= {16'd72, 16'd32767};
                15'd24 : data_rom <= {16'd75, 16'd32767};
                15'd25 : data_rom <= {16'd78, 16'd32767};
                15'd26 : data_rom <= {16'd81, 16'd32767};
                15'd27 : data_rom <= {16'd84, 16'd32767};
                15'd28 : data_rom <= {16'd87, 16'd32767};
                15'd29 : data_rom <= {16'd91, 16'd32767};
                15'd30 : data_rom <= {16'd94, 16'd32767};
                15'd31 : data_rom <= {16'd97, 16'd32767};
                15'd32 : data_rom <= {16'd100, 16'd32767};
                15'd33 : data_rom <= {16'd103, 16'd32767};
                15'd34 : data_rom <= {16'd106, 16'd32767};
                15'd35 : data_rom <= {16'd109, 16'd32767};
                15'd36 : data_rom <= {16'd113, 16'd32767};
                15'd37 : data_rom <= {16'd116, 16'd32767};
                15'd38 : data_rom <= {16'd119, 16'd32767};
                15'd39 : data_rom <= {16'd122, 16'd32767};
                15'd40 : data_rom <= {16'd125, 16'd32767};
                15'd41 : data_rom <= {16'd128, 16'd32767};
                15'd42 : data_rom <= {16'd131, 16'd32767};
                15'd43 : data_rom <= {16'd135, 16'd32767};
                15'd44 : data_rom <= {16'd138, 16'd32767};
                15'd45 : data_rom <= {16'd141, 16'd32767};
                15'd46 : data_rom <= {16'd144, 16'd32767};
                15'd47 : data_rom <= {16'd147, 16'd32767};
                15'd48 : data_rom <= {16'd150, 16'd32767};
                15'd49 : data_rom <= {16'd153, 16'd32767};
                15'd50 : data_rom <= {16'd157, 16'd32767};
                15'd51 : data_rom <= {16'd160, 16'd32767};
                15'd52 : data_rom <= {16'd163, 16'd32767};
                15'd53 : data_rom <= {16'd166, 16'd32767};
                15'd54 : data_rom <= {16'd169, 16'd32767};
                15'd55 : data_rom <= {16'd172, 16'd32767};
                15'd56 : data_rom <= {16'd175, 16'd32767};
                15'd57 : data_rom <= {16'd179, 16'd32767};
                15'd58 : data_rom <= {16'd182, 16'd32767};
                15'd59 : data_rom <= {16'd185, 16'd32767};
                15'd60 : data_rom <= {16'd188, 16'd32767};
                15'd61 : data_rom <= {16'd191, 16'd32767};
                15'd62 : data_rom <= {16'd194, 16'd32767};
                15'd63 : data_rom <= {16'd197, 16'd32767};
                15'd64 : data_rom <= {16'd201, 16'd32767};
                15'd65 : data_rom <= {16'd204, 16'd32767};
                15'd66 : data_rom <= {16'd207, 16'd32767};
                15'd67 : data_rom <= {16'd210, 16'd32767};
                15'd68 : data_rom <= {16'd213, 16'd32767};
                15'd69 : data_rom <= {16'd216, 16'd32767};
                15'd70 : data_rom <= {16'd219, 16'd32767};
                15'd71 : data_rom <= {16'd223, 16'd32767};
                15'd72 : data_rom <= {16'd226, 16'd32767};
                15'd73 : data_rom <= {16'd229, 16'd32767};
                15'd74 : data_rom <= {16'd232, 16'd32767};
                15'd75 : data_rom <= {16'd235, 16'd32767};
                15'd76 : data_rom <= {16'd238, 16'd32767};
                15'd77 : data_rom <= {16'd241, 16'd32767};
                15'd78 : data_rom <= {16'd245, 16'd32767};
                15'd79 : data_rom <= {16'd248, 16'd32767};
                15'd80 : data_rom <= {16'd251, 16'd32767};
                15'd81 : data_rom <= {16'd254, 16'd32767};
                15'd82 : data_rom <= {16'd257, 16'd32766};
                15'd83 : data_rom <= {16'd260, 16'd32766};
                15'd84 : data_rom <= {16'd263, 16'd32766};
                15'd85 : data_rom <= {16'd267, 16'd32766};
                15'd86 : data_rom <= {16'd270, 16'd32766};
                15'd87 : data_rom <= {16'd273, 16'd32766};
                15'd88 : data_rom <= {16'd276, 16'd32766};
                15'd89 : data_rom <= {16'd279, 16'd32766};
                15'd90 : data_rom <= {16'd282, 16'd32766};
                15'd91 : data_rom <= {16'd285, 16'd32766};
                15'd92 : data_rom <= {16'd289, 16'd32766};
                15'd93 : data_rom <= {16'd292, 16'd32766};
                15'd94 : data_rom <= {16'd295, 16'd32766};
                15'd95 : data_rom <= {16'd298, 16'd32766};
                15'd96 : data_rom <= {16'd301, 16'd32766};
                15'd97 : data_rom <= {16'd304, 16'd32766};
                15'd98 : data_rom <= {16'd307, 16'd32766};
                15'd99 : data_rom <= {16'd311, 16'd32766};
                15'd100 : data_rom <= {16'd314, 16'd32766};
                15'd101 : data_rom <= {16'd317, 16'd32766};
                15'd102 : data_rom <= {16'd320, 16'd32766};
                15'd103 : data_rom <= {16'd323, 16'd32766};
                15'd104 : data_rom <= {16'd326, 16'd32766};
                15'd105 : data_rom <= {16'd329, 16'd32766};
                15'd106 : data_rom <= {16'd333, 16'd32766};
                15'd107 : data_rom <= {16'd336, 16'd32766};
                15'd108 : data_rom <= {16'd339, 16'd32766};
                15'd109 : data_rom <= {16'd342, 16'd32766};
                15'd110 : data_rom <= {16'd345, 16'd32766};
                15'd111 : data_rom <= {16'd348, 16'd32766};
                15'd112 : data_rom <= {16'd351, 16'd32766};
                15'd113 : data_rom <= {16'd354, 16'd32766};
                15'd114 : data_rom <= {16'd358, 16'd32766};
                15'd115 : data_rom <= {16'd361, 16'd32766};
                15'd116 : data_rom <= {16'd364, 16'd32765};
                15'd117 : data_rom <= {16'd367, 16'd32765};
                15'd118 : data_rom <= {16'd370, 16'd32765};
                15'd119 : data_rom <= {16'd373, 16'd32765};
                15'd120 : data_rom <= {16'd376, 16'd32765};
                15'd121 : data_rom <= {16'd380, 16'd32765};
                15'd122 : data_rom <= {16'd383, 16'd32765};
                15'd123 : data_rom <= {16'd386, 16'd32765};
                15'd124 : data_rom <= {16'd389, 16'd32765};
                15'd125 : data_rom <= {16'd392, 16'd32765};
                15'd126 : data_rom <= {16'd395, 16'd32765};
                15'd127 : data_rom <= {16'd398, 16'd32765};
                15'd128 : data_rom <= {16'd402, 16'd32765};
                15'd129 : data_rom <= {16'd405, 16'd32765};
                15'd130 : data_rom <= {16'd408, 16'd32765};
                15'd131 : data_rom <= {16'd411, 16'd32765};
                15'd132 : data_rom <= {16'd414, 16'd32765};
                15'd133 : data_rom <= {16'd417, 16'd32765};
                15'd134 : data_rom <= {16'd420, 16'd32765};
                15'd135 : data_rom <= {16'd424, 16'd32765};
                15'd136 : data_rom <= {16'd427, 16'd32765};
                15'd137 : data_rom <= {16'd430, 16'd32765};
                15'd138 : data_rom <= {16'd433, 16'd32765};
                15'd139 : data_rom <= {16'd436, 16'd32765};
                15'd140 : data_rom <= {16'd439, 16'd32765};
                15'd141 : data_rom <= {16'd442, 16'd32765};
                15'd142 : data_rom <= {16'd446, 16'd32764};
                15'd143 : data_rom <= {16'd449, 16'd32764};
                15'd144 : data_rom <= {16'd452, 16'd32764};
                15'd145 : data_rom <= {16'd455, 16'd32764};
                15'd146 : data_rom <= {16'd458, 16'd32764};
                15'd147 : data_rom <= {16'd461, 16'd32764};
                15'd148 : data_rom <= {16'd464, 16'd32764};
                15'd149 : data_rom <= {16'd468, 16'd32764};
                15'd150 : data_rom <= {16'd471, 16'd32764};
                15'd151 : data_rom <= {16'd474, 16'd32764};
                15'd152 : data_rom <= {16'd477, 16'd32764};
                15'd153 : data_rom <= {16'd480, 16'd32764};
                15'd154 : data_rom <= {16'd483, 16'd32764};
                15'd155 : data_rom <= {16'd486, 16'd32764};
                15'd156 : data_rom <= {16'd490, 16'd32764};
                15'd157 : data_rom <= {16'd493, 16'd32764};
                15'd158 : data_rom <= {16'd496, 16'd32764};
                15'd159 : data_rom <= {16'd499, 16'd32764};
                15'd160 : data_rom <= {16'd502, 16'd32764};
                15'd161 : data_rom <= {16'd505, 16'd32764};
                15'd162 : data_rom <= {16'd508, 16'd32764};
                15'd163 : data_rom <= {16'd512, 16'd32763};
                15'd164 : data_rom <= {16'd515, 16'd32763};
                15'd165 : data_rom <= {16'd518, 16'd32763};
                15'd166 : data_rom <= {16'd521, 16'd32763};
                15'd167 : data_rom <= {16'd524, 16'd32763};
                15'd168 : data_rom <= {16'd527, 16'd32763};
                15'd169 : data_rom <= {16'd530, 16'd32763};
                15'd170 : data_rom <= {16'd534, 16'd32763};
                15'd171 : data_rom <= {16'd537, 16'd32763};
                15'd172 : data_rom <= {16'd540, 16'd32763};
                15'd173 : data_rom <= {16'd543, 16'd32763};
                15'd174 : data_rom <= {16'd546, 16'd32763};
                15'd175 : data_rom <= {16'd549, 16'd32763};
                15'd176 : data_rom <= {16'd552, 16'd32763};
                15'd177 : data_rom <= {16'd556, 16'd32763};
                15'd178 : data_rom <= {16'd559, 16'd32763};
                15'd179 : data_rom <= {16'd562, 16'd32763};
                15'd180 : data_rom <= {16'd565, 16'd32763};
                15'd181 : data_rom <= {16'd568, 16'd32763};
                15'd182 : data_rom <= {16'd571, 16'd32763};
                15'd183 : data_rom <= {16'd574, 16'd32762};
                15'd184 : data_rom <= {16'd578, 16'd32762};
                15'd185 : data_rom <= {16'd581, 16'd32762};
                15'd186 : data_rom <= {16'd584, 16'd32762};
                15'd187 : data_rom <= {16'd587, 16'd32762};
                15'd188 : data_rom <= {16'd590, 16'd32762};
                15'd189 : data_rom <= {16'd593, 16'd32762};
                15'd190 : data_rom <= {16'd596, 16'd32762};
                15'd191 : data_rom <= {16'd600, 16'd32762};
                15'd192 : data_rom <= {16'd603, 16'd32762};
                15'd193 : data_rom <= {16'd606, 16'd32762};
                15'd194 : data_rom <= {16'd609, 16'd32762};
                15'd195 : data_rom <= {16'd612, 16'd32762};
                15'd196 : data_rom <= {16'd615, 16'd32762};
                15'd197 : data_rom <= {16'd618, 16'd32762};
                15'd198 : data_rom <= {16'd621, 16'd32762};
                15'd199 : data_rom <= {16'd625, 16'd32762};
                15'd200 : data_rom <= {16'd628, 16'd32761};
                15'd201 : data_rom <= {16'd631, 16'd32761};
                15'd202 : data_rom <= {16'd634, 16'd32761};
                15'd203 : data_rom <= {16'd637, 16'd32761};
                15'd204 : data_rom <= {16'd640, 16'd32761};
                15'd205 : data_rom <= {16'd643, 16'd32761};
                15'd206 : data_rom <= {16'd647, 16'd32761};
                15'd207 : data_rom <= {16'd650, 16'd32761};
                15'd208 : data_rom <= {16'd653, 16'd32761};
                15'd209 : data_rom <= {16'd656, 16'd32761};
                15'd210 : data_rom <= {16'd659, 16'd32761};
                15'd211 : data_rom <= {16'd662, 16'd32761};
                15'd212 : data_rom <= {16'd665, 16'd32761};
                15'd213 : data_rom <= {16'd669, 16'd32761};
                15'd214 : data_rom <= {16'd672, 16'd32761};
                15'd215 : data_rom <= {16'd675, 16'd32761};
                15'd216 : data_rom <= {16'd678, 16'd32760};
                15'd217 : data_rom <= {16'd681, 16'd32760};
                15'd218 : data_rom <= {16'd684, 16'd32760};
                15'd219 : data_rom <= {16'd687, 16'd32760};
                15'd220 : data_rom <= {16'd691, 16'd32760};
                15'd221 : data_rom <= {16'd694, 16'd32760};
                15'd222 : data_rom <= {16'd697, 16'd32760};
                15'd223 : data_rom <= {16'd700, 16'd32760};
                15'd224 : data_rom <= {16'd703, 16'd32760};
                15'd225 : data_rom <= {16'd706, 16'd32760};
                15'd226 : data_rom <= {16'd709, 16'd32760};
                15'd227 : data_rom <= {16'd713, 16'd32760};
                15'd228 : data_rom <= {16'd716, 16'd32760};
                15'd229 : data_rom <= {16'd719, 16'd32760};
                15'd230 : data_rom <= {16'd722, 16'd32760};
                15'd231 : data_rom <= {16'd725, 16'd32759};
                15'd232 : data_rom <= {16'd728, 16'd32759};
                15'd233 : data_rom <= {16'd731, 16'd32759};
                15'd234 : data_rom <= {16'd735, 16'd32759};
                15'd235 : data_rom <= {16'd738, 16'd32759};
                15'd236 : data_rom <= {16'd741, 16'd32759};
                15'd237 : data_rom <= {16'd744, 16'd32759};
                15'd238 : data_rom <= {16'd747, 16'd32759};
                15'd239 : data_rom <= {16'd750, 16'd32759};
                15'd240 : data_rom <= {16'd753, 16'd32759};
                15'd241 : data_rom <= {16'd757, 16'd32759};
                15'd242 : data_rom <= {16'd760, 16'd32759};
                15'd243 : data_rom <= {16'd763, 16'd32759};
                15'd244 : data_rom <= {16'd766, 16'd32759};
                15'd245 : data_rom <= {16'd769, 16'd32758};
                15'd246 : data_rom <= {16'd772, 16'd32758};
                15'd247 : data_rom <= {16'd775, 16'd32758};
                15'd248 : data_rom <= {16'd779, 16'd32758};
                15'd249 : data_rom <= {16'd782, 16'd32758};
                15'd250 : data_rom <= {16'd785, 16'd32758};
                15'd251 : data_rom <= {16'd788, 16'd32758};
                15'd252 : data_rom <= {16'd791, 16'd32758};
                15'd253 : data_rom <= {16'd794, 16'd32758};
                15'd254 : data_rom <= {16'd797, 16'd32758};
                15'd255 : data_rom <= {16'd801, 16'd32758};
                15'd256 : data_rom <= {16'd804, 16'd32758};
                15'd257 : data_rom <= {16'd807, 16'd32758};
                15'd258 : data_rom <= {16'd810, 16'd32757};
                15'd259 : data_rom <= {16'd813, 16'd32757};
                15'd260 : data_rom <= {16'd816, 16'd32757};
                15'd261 : data_rom <= {16'd819, 16'd32757};
                15'd262 : data_rom <= {16'd823, 16'd32757};
                15'd263 : data_rom <= {16'd826, 16'd32757};
                15'd264 : data_rom <= {16'd829, 16'd32757};
                15'd265 : data_rom <= {16'd832, 16'd32757};
                15'd266 : data_rom <= {16'd835, 16'd32757};
                15'd267 : data_rom <= {16'd838, 16'd32757};
                15'd268 : data_rom <= {16'd841, 16'd32757};
                15'd269 : data_rom <= {16'd844, 16'd32757};
                15'd270 : data_rom <= {16'd848, 16'd32757};
                15'd271 : data_rom <= {16'd851, 16'd32756};
                15'd272 : data_rom <= {16'd854, 16'd32756};
                15'd273 : data_rom <= {16'd857, 16'd32756};
                15'd274 : data_rom <= {16'd860, 16'd32756};
                15'd275 : data_rom <= {16'd863, 16'd32756};
                15'd276 : data_rom <= {16'd866, 16'd32756};
                15'd277 : data_rom <= {16'd870, 16'd32756};
                15'd278 : data_rom <= {16'd873, 16'd32756};
                15'd279 : data_rom <= {16'd876, 16'd32756};
                15'd280 : data_rom <= {16'd879, 16'd32756};
                15'd281 : data_rom <= {16'd882, 16'd32756};
                15'd282 : data_rom <= {16'd885, 16'd32756};
                15'd283 : data_rom <= {16'd888, 16'd32755};
                15'd284 : data_rom <= {16'd892, 16'd32755};
                15'd285 : data_rom <= {16'd895, 16'd32755};
                15'd286 : data_rom <= {16'd898, 16'd32755};
                15'd287 : data_rom <= {16'd901, 16'd32755};
                15'd288 : data_rom <= {16'd904, 16'd32755};
                15'd289 : data_rom <= {16'd907, 16'd32755};
                15'd290 : data_rom <= {16'd910, 16'd32755};
                15'd291 : data_rom <= {16'd914, 16'd32755};
                15'd292 : data_rom <= {16'd917, 16'd32755};
                15'd293 : data_rom <= {16'd920, 16'd32755};
                15'd294 : data_rom <= {16'd923, 16'd32754};
                15'd295 : data_rom <= {16'd926, 16'd32754};
                15'd296 : data_rom <= {16'd929, 16'd32754};
                15'd297 : data_rom <= {16'd932, 16'd32754};
                15'd298 : data_rom <= {16'd936, 16'd32754};
                15'd299 : data_rom <= {16'd939, 16'd32754};
                15'd300 : data_rom <= {16'd942, 16'd32754};
                15'd301 : data_rom <= {16'd945, 16'd32754};
                15'd302 : data_rom <= {16'd948, 16'd32754};
                15'd303 : data_rom <= {16'd951, 16'd32754};
                15'd304 : data_rom <= {16'd954, 16'd32754};
                15'd305 : data_rom <= {16'd958, 16'd32753};
                15'd306 : data_rom <= {16'd961, 16'd32753};
                15'd307 : data_rom <= {16'd964, 16'd32753};
                15'd308 : data_rom <= {16'd967, 16'd32753};
                15'd309 : data_rom <= {16'd970, 16'd32753};
                15'd310 : data_rom <= {16'd973, 16'd32753};
                15'd311 : data_rom <= {16'd976, 16'd32753};
                15'd312 : data_rom <= {16'd980, 16'd32753};
                15'd313 : data_rom <= {16'd983, 16'd32753};
                15'd314 : data_rom <= {16'd986, 16'd32753};
                15'd315 : data_rom <= {16'd989, 16'd32753};
                15'd316 : data_rom <= {16'd992, 16'd32752};
                15'd317 : data_rom <= {16'd995, 16'd32752};
                15'd318 : data_rom <= {16'd998, 16'd32752};
                15'd319 : data_rom <= {16'd1002, 16'd32752};
                15'd320 : data_rom <= {16'd1005, 16'd32752};
                15'd321 : data_rom <= {16'd1008, 16'd32752};
                15'd322 : data_rom <= {16'd1011, 16'd32752};
                15'd323 : data_rom <= {16'd1014, 16'd32752};
                15'd324 : data_rom <= {16'd1017, 16'd32752};
                15'd325 : data_rom <= {16'd1020, 16'd32752};
                15'd326 : data_rom <= {16'd1023, 16'd32751};
                15'd327 : data_rom <= {16'd1027, 16'd32751};
                15'd328 : data_rom <= {16'd1030, 16'd32751};
                15'd329 : data_rom <= {16'd1033, 16'd32751};
                15'd330 : data_rom <= {16'd1036, 16'd32751};
                15'd331 : data_rom <= {16'd1039, 16'd32751};
                15'd332 : data_rom <= {16'd1042, 16'd32751};
                15'd333 : data_rom <= {16'd1045, 16'd32751};
                15'd334 : data_rom <= {16'd1049, 16'd32751};
                15'd335 : data_rom <= {16'd1052, 16'd32751};
                15'd336 : data_rom <= {16'd1055, 16'd32750};
                15'd337 : data_rom <= {16'd1058, 16'd32750};
                15'd338 : data_rom <= {16'd1061, 16'd32750};
                15'd339 : data_rom <= {16'd1064, 16'd32750};
                15'd340 : data_rom <= {16'd1067, 16'd32750};
                15'd341 : data_rom <= {16'd1071, 16'd32750};
                15'd342 : data_rom <= {16'd1074, 16'd32750};
                15'd343 : data_rom <= {16'd1077, 16'd32750};
                15'd344 : data_rom <= {16'd1080, 16'd32750};
                15'd345 : data_rom <= {16'd1083, 16'd32750};
                15'd346 : data_rom <= {16'd1086, 16'd32749};
                15'd347 : data_rom <= {16'd1089, 16'd32749};
                15'd348 : data_rom <= {16'd1093, 16'd32749};
                15'd349 : data_rom <= {16'd1096, 16'd32749};
                15'd350 : data_rom <= {16'd1099, 16'd32749};
                15'd351 : data_rom <= {16'd1102, 16'd32749};
                15'd352 : data_rom <= {16'd1105, 16'd32749};
                15'd353 : data_rom <= {16'd1108, 16'd32749};
                15'd354 : data_rom <= {16'd1111, 16'd32749};
                15'd355 : data_rom <= {16'd1115, 16'd32749};
                15'd356 : data_rom <= {16'd1118, 16'd32748};
                15'd357 : data_rom <= {16'd1121, 16'd32748};
                15'd358 : data_rom <= {16'd1124, 16'd32748};
                15'd359 : data_rom <= {16'd1127, 16'd32748};
                15'd360 : data_rom <= {16'd1130, 16'd32748};
                15'd361 : data_rom <= {16'd1133, 16'd32748};
                15'd362 : data_rom <= {16'd1137, 16'd32748};
                15'd363 : data_rom <= {16'd1140, 16'd32748};
                15'd364 : data_rom <= {16'd1143, 16'd32748};
                15'd365 : data_rom <= {16'd1146, 16'd32747};
                15'd366 : data_rom <= {16'd1149, 16'd32747};
                15'd367 : data_rom <= {16'd1152, 16'd32747};
                15'd368 : data_rom <= {16'd1155, 16'd32747};
                15'd369 : data_rom <= {16'd1159, 16'd32747};
                15'd370 : data_rom <= {16'd1162, 16'd32747};
                15'd371 : data_rom <= {16'd1165, 16'd32747};
                15'd372 : data_rom <= {16'd1168, 16'd32747};
                15'd373 : data_rom <= {16'd1171, 16'd32747};
                15'd374 : data_rom <= {16'd1174, 16'd32746};
                15'd375 : data_rom <= {16'd1177, 16'd32746};
                15'd376 : data_rom <= {16'd1180, 16'd32746};
                15'd377 : data_rom <= {16'd1184, 16'd32746};
                15'd378 : data_rom <= {16'd1187, 16'd32746};
                15'd379 : data_rom <= {16'd1190, 16'd32746};
                15'd380 : data_rom <= {16'd1193, 16'd32746};
                15'd381 : data_rom <= {16'd1196, 16'd32746};
                15'd382 : data_rom <= {16'd1199, 16'd32746};
                15'd383 : data_rom <= {16'd1202, 16'd32745};
                15'd384 : data_rom <= {16'd1206, 16'd32745};
                15'd385 : data_rom <= {16'd1209, 16'd32745};
                15'd386 : data_rom <= {16'd1212, 16'd32745};
                15'd387 : data_rom <= {16'd1215, 16'd32745};
                15'd388 : data_rom <= {16'd1218, 16'd32745};
                15'd389 : data_rom <= {16'd1221, 16'd32745};
                15'd390 : data_rom <= {16'd1224, 16'd32745};
                15'd391 : data_rom <= {16'd1228, 16'd32744};
                15'd392 : data_rom <= {16'd1231, 16'd32744};
                15'd393 : data_rom <= {16'd1234, 16'd32744};
                15'd394 : data_rom <= {16'd1237, 16'd32744};
                15'd395 : data_rom <= {16'd1240, 16'd32744};
                15'd396 : data_rom <= {16'd1243, 16'd32744};
                15'd397 : data_rom <= {16'd1246, 16'd32744};
                15'd398 : data_rom <= {16'd1250, 16'd32744};
                15'd399 : data_rom <= {16'd1253, 16'd32744};
                15'd400 : data_rom <= {16'd1256, 16'd32743};
                15'd401 : data_rom <= {16'd1259, 16'd32743};
                15'd402 : data_rom <= {16'd1262, 16'd32743};
                15'd403 : data_rom <= {16'd1265, 16'd32743};
                15'd404 : data_rom <= {16'd1268, 16'd32743};
                15'd405 : data_rom <= {16'd1272, 16'd32743};
                15'd406 : data_rom <= {16'd1275, 16'd32743};
                15'd407 : data_rom <= {16'd1278, 16'd32743};
                15'd408 : data_rom <= {16'd1281, 16'd32742};
                15'd409 : data_rom <= {16'd1284, 16'd32742};
                15'd410 : data_rom <= {16'd1287, 16'd32742};
                15'd411 : data_rom <= {16'd1290, 16'd32742};
                15'd412 : data_rom <= {16'd1293, 16'd32742};
                15'd413 : data_rom <= {16'd1297, 16'd32742};
                15'd414 : data_rom <= {16'd1300, 16'd32742};
                15'd415 : data_rom <= {16'd1303, 16'd32742};
                15'd416 : data_rom <= {16'd1306, 16'd32741};
                15'd417 : data_rom <= {16'd1309, 16'd32741};
                15'd418 : data_rom <= {16'd1312, 16'd32741};
                15'd419 : data_rom <= {16'd1315, 16'd32741};
                15'd420 : data_rom <= {16'd1319, 16'd32741};
                15'd421 : data_rom <= {16'd1322, 16'd32741};
                15'd422 : data_rom <= {16'd1325, 16'd32741};
                15'd423 : data_rom <= {16'd1328, 16'd32741};
                15'd424 : data_rom <= {16'd1331, 16'd32740};
                15'd425 : data_rom <= {16'd1334, 16'd32740};
                15'd426 : data_rom <= {16'd1337, 16'd32740};
                15'd427 : data_rom <= {16'd1341, 16'd32740};
                15'd428 : data_rom <= {16'd1344, 16'd32740};
                15'd429 : data_rom <= {16'd1347, 16'd32740};
                15'd430 : data_rom <= {16'd1350, 16'd32740};
                15'd431 : data_rom <= {16'd1353, 16'd32740};
                15'd432 : data_rom <= {16'd1356, 16'd32739};
                15'd433 : data_rom <= {16'd1359, 16'd32739};
                15'd434 : data_rom <= {16'd1363, 16'd32739};
                15'd435 : data_rom <= {16'd1366, 16'd32739};
                15'd436 : data_rom <= {16'd1369, 16'd32739};
                15'd437 : data_rom <= {16'd1372, 16'd32739};
                15'd438 : data_rom <= {16'd1375, 16'd32739};
                15'd439 : data_rom <= {16'd1378, 16'd32738};
                15'd440 : data_rom <= {16'd1381, 16'd32738};
                15'd441 : data_rom <= {16'd1385, 16'd32738};
                15'd442 : data_rom <= {16'd1388, 16'd32738};
                15'd443 : data_rom <= {16'd1391, 16'd32738};
                15'd444 : data_rom <= {16'd1394, 16'd32738};
                15'd445 : data_rom <= {16'd1397, 16'd32738};
                15'd446 : data_rom <= {16'd1400, 16'd32738};
                15'd447 : data_rom <= {16'd1403, 16'd32737};
                15'd448 : data_rom <= {16'd1406, 16'd32737};
                15'd449 : data_rom <= {16'd1410, 16'd32737};
                15'd450 : data_rom <= {16'd1413, 16'd32737};
                15'd451 : data_rom <= {16'd1416, 16'd32737};
                15'd452 : data_rom <= {16'd1419, 16'd32737};
                15'd453 : data_rom <= {16'd1422, 16'd32737};
                15'd454 : data_rom <= {16'd1425, 16'd32736};
                15'd455 : data_rom <= {16'd1428, 16'd32736};
                15'd456 : data_rom <= {16'd1432, 16'd32736};
                15'd457 : data_rom <= {16'd1435, 16'd32736};
                15'd458 : data_rom <= {16'd1438, 16'd32736};
                15'd459 : data_rom <= {16'd1441, 16'd32736};
                15'd460 : data_rom <= {16'd1444, 16'd32736};
                15'd461 : data_rom <= {16'd1447, 16'd32735};
                15'd462 : data_rom <= {16'd1450, 16'd32735};
                15'd463 : data_rom <= {16'd1454, 16'd32735};
                15'd464 : data_rom <= {16'd1457, 16'd32735};
                15'd465 : data_rom <= {16'd1460, 16'd32735};
                15'd466 : data_rom <= {16'd1463, 16'd32735};
                15'd467 : data_rom <= {16'd1466, 16'd32735};
                15'd468 : data_rom <= {16'd1469, 16'd32735};
                15'd469 : data_rom <= {16'd1472, 16'd32734};
                15'd470 : data_rom <= {16'd1476, 16'd32734};
                15'd471 : data_rom <= {16'd1479, 16'd32734};
                15'd472 : data_rom <= {16'd1482, 16'd32734};
                15'd473 : data_rom <= {16'd1485, 16'd32734};
                15'd474 : data_rom <= {16'd1488, 16'd32734};
                15'd475 : data_rom <= {16'd1491, 16'd32734};
                15'd476 : data_rom <= {16'd1494, 16'd32733};
                15'd477 : data_rom <= {16'd1498, 16'd32733};
                15'd478 : data_rom <= {16'd1501, 16'd32733};
                15'd479 : data_rom <= {16'd1504, 16'd32733};
                15'd480 : data_rom <= {16'd1507, 16'd32733};
                15'd481 : data_rom <= {16'd1510, 16'd32733};
                15'd482 : data_rom <= {16'd1513, 16'd32733};
                15'd483 : data_rom <= {16'd1516, 16'd32732};
                15'd484 : data_rom <= {16'd1519, 16'd32732};
                15'd485 : data_rom <= {16'd1523, 16'd32732};
                15'd486 : data_rom <= {16'd1526, 16'd32732};
                15'd487 : data_rom <= {16'd1529, 16'd32732};
                15'd488 : data_rom <= {16'd1532, 16'd32732};
                15'd489 : data_rom <= {16'd1535, 16'd32731};
                15'd490 : data_rom <= {16'd1538, 16'd32731};
                15'd491 : data_rom <= {16'd1541, 16'd32731};
                15'd492 : data_rom <= {16'd1545, 16'd32731};
                15'd493 : data_rom <= {16'd1548, 16'd32731};
                15'd494 : data_rom <= {16'd1551, 16'd32731};
                15'd495 : data_rom <= {16'd1554, 16'd32731};
                15'd496 : data_rom <= {16'd1557, 16'd32730};
                15'd497 : data_rom <= {16'd1560, 16'd32730};
                15'd498 : data_rom <= {16'd1563, 16'd32730};
                15'd499 : data_rom <= {16'd1567, 16'd32730};
                15'd500 : data_rom <= {16'd1570, 16'd32730};
                15'd501 : data_rom <= {16'd1573, 16'd32730};
                15'd502 : data_rom <= {16'd1576, 16'd32730};
                15'd503 : data_rom <= {16'd1579, 16'd32729};
                15'd504 : data_rom <= {16'd1582, 16'd32729};
                15'd505 : data_rom <= {16'd1585, 16'd32729};
                15'd506 : data_rom <= {16'd1589, 16'd32729};
                15'd507 : data_rom <= {16'd1592, 16'd32729};
                15'd508 : data_rom <= {16'd1595, 16'd32729};
                15'd509 : data_rom <= {16'd1598, 16'd32728};
                15'd510 : data_rom <= {16'd1601, 16'd32728};
                15'd511 : data_rom <= {16'd1604, 16'd32728};
                15'd512 : data_rom <= {16'd1607, 16'd32728};
                15'd513 : data_rom <= {16'd1610, 16'd32728};
                15'd514 : data_rom <= {16'd1614, 16'd32728};
                15'd515 : data_rom <= {16'd1617, 16'd32728};
                15'd516 : data_rom <= {16'd1620, 16'd32727};
                15'd517 : data_rom <= {16'd1623, 16'd32727};
                15'd518 : data_rom <= {16'd1626, 16'd32727};
                15'd519 : data_rom <= {16'd1629, 16'd32727};
                15'd520 : data_rom <= {16'd1632, 16'd32727};
                15'd521 : data_rom <= {16'd1636, 16'd32727};
                15'd522 : data_rom <= {16'd1639, 16'd32726};
                15'd523 : data_rom <= {16'd1642, 16'd32726};
                15'd524 : data_rom <= {16'd1645, 16'd32726};
                15'd525 : data_rom <= {16'd1648, 16'd32726};
                15'd526 : data_rom <= {16'd1651, 16'd32726};
                15'd527 : data_rom <= {16'd1654, 16'd32726};
                15'd528 : data_rom <= {16'd1658, 16'd32726};
                15'd529 : data_rom <= {16'd1661, 16'd32725};
                15'd530 : data_rom <= {16'd1664, 16'd32725};
                15'd531 : data_rom <= {16'd1667, 16'd32725};
                15'd532 : data_rom <= {16'd1670, 16'd32725};
                15'd533 : data_rom <= {16'd1673, 16'd32725};
                15'd534 : data_rom <= {16'd1676, 16'd32725};
                15'd535 : data_rom <= {16'd1680, 16'd32724};
                15'd536 : data_rom <= {16'd1683, 16'd32724};
                15'd537 : data_rom <= {16'd1686, 16'd32724};
                15'd538 : data_rom <= {16'd1689, 16'd32724};
                15'd539 : data_rom <= {16'd1692, 16'd32724};
                15'd540 : data_rom <= {16'd1695, 16'd32724};
                15'd541 : data_rom <= {16'd1698, 16'd32723};
                15'd542 : data_rom <= {16'd1701, 16'd32723};
                15'd543 : data_rom <= {16'd1705, 16'd32723};
                15'd544 : data_rom <= {16'd1708, 16'd32723};
                15'd545 : data_rom <= {16'd1711, 16'd32723};
                15'd546 : data_rom <= {16'd1714, 16'd32723};
                15'd547 : data_rom <= {16'd1717, 16'd32722};
                15'd548 : data_rom <= {16'd1720, 16'd32722};
                15'd549 : data_rom <= {16'd1723, 16'd32722};
                15'd550 : data_rom <= {16'd1727, 16'd32722};
                15'd551 : data_rom <= {16'd1730, 16'd32722};
                15'd552 : data_rom <= {16'd1733, 16'd32722};
                15'd553 : data_rom <= {16'd1736, 16'd32721};
                15'd554 : data_rom <= {16'd1739, 16'd32721};
                15'd555 : data_rom <= {16'd1742, 16'd32721};
                15'd556 : data_rom <= {16'd1745, 16'd32721};
                15'd557 : data_rom <= {16'd1749, 16'd32721};
                15'd558 : data_rom <= {16'd1752, 16'd32721};
                15'd559 : data_rom <= {16'd1755, 16'd32720};
                15'd560 : data_rom <= {16'd1758, 16'd32720};
                15'd561 : data_rom <= {16'd1761, 16'd32720};
                15'd562 : data_rom <= {16'd1764, 16'd32720};
                15'd563 : data_rom <= {16'd1767, 16'd32720};
                15'd564 : data_rom <= {16'd1770, 16'd32720};
                15'd565 : data_rom <= {16'd1774, 16'd32719};
                15'd566 : data_rom <= {16'd1777, 16'd32719};
                15'd567 : data_rom <= {16'd1780, 16'd32719};
                15'd568 : data_rom <= {16'd1783, 16'd32719};
                15'd569 : data_rom <= {16'd1786, 16'd32719};
                15'd570 : data_rom <= {16'd1789, 16'd32719};
                15'd571 : data_rom <= {16'd1792, 16'd32718};
                15'd572 : data_rom <= {16'd1796, 16'd32718};
                15'd573 : data_rom <= {16'd1799, 16'd32718};
                15'd574 : data_rom <= {16'd1802, 16'd32718};
                15'd575 : data_rom <= {16'd1805, 16'd32718};
                15'd576 : data_rom <= {16'd1808, 16'd32718};
                15'd577 : data_rom <= {16'd1811, 16'd32717};
                15'd578 : data_rom <= {16'd1814, 16'd32717};
                15'd579 : data_rom <= {16'd1818, 16'd32717};
                15'd580 : data_rom <= {16'd1821, 16'd32717};
                15'd581 : data_rom <= {16'd1824, 16'd32717};
                15'd582 : data_rom <= {16'd1827, 16'd32717};
                15'd583 : data_rom <= {16'd1830, 16'd32716};
                15'd584 : data_rom <= {16'd1833, 16'd32716};
                15'd585 : data_rom <= {16'd1836, 16'd32716};
                15'd586 : data_rom <= {16'd1840, 16'd32716};
                15'd587 : data_rom <= {16'd1843, 16'd32716};
                15'd588 : data_rom <= {16'd1846, 16'd32715};
                15'd589 : data_rom <= {16'd1849, 16'd32715};
                15'd590 : data_rom <= {16'd1852, 16'd32715};
                15'd591 : data_rom <= {16'd1855, 16'd32715};
                15'd592 : data_rom <= {16'd1858, 16'd32715};
                15'd593 : data_rom <= {16'd1861, 16'd32715};
                15'd594 : data_rom <= {16'd1865, 16'd32714};
                15'd595 : data_rom <= {16'd1868, 16'd32714};
                15'd596 : data_rom <= {16'd1871, 16'd32714};
                15'd597 : data_rom <= {16'd1874, 16'd32714};
                15'd598 : data_rom <= {16'd1877, 16'd32714};
                15'd599 : data_rom <= {16'd1880, 16'd32713};
                15'd600 : data_rom <= {16'd1883, 16'd32713};
                15'd601 : data_rom <= {16'd1887, 16'd32713};
                15'd602 : data_rom <= {16'd1890, 16'd32713};
                15'd603 : data_rom <= {16'd1893, 16'd32713};
                15'd604 : data_rom <= {16'd1896, 16'd32713};
                15'd605 : data_rom <= {16'd1899, 16'd32712};
                15'd606 : data_rom <= {16'd1902, 16'd32712};
                15'd607 : data_rom <= {16'd1905, 16'd32712};
                15'd608 : data_rom <= {16'd1909, 16'd32712};
                15'd609 : data_rom <= {16'd1912, 16'd32712};
                15'd610 : data_rom <= {16'd1915, 16'd32711};
                15'd611 : data_rom <= {16'd1918, 16'd32711};
                15'd612 : data_rom <= {16'd1921, 16'd32711};
                15'd613 : data_rom <= {16'd1924, 16'd32711};
                15'd614 : data_rom <= {16'd1927, 16'd32711};
                15'd615 : data_rom <= {16'd1930, 16'd32711};
                15'd616 : data_rom <= {16'd1934, 16'd32710};
                15'd617 : data_rom <= {16'd1937, 16'd32710};
                15'd618 : data_rom <= {16'd1940, 16'd32710};
                15'd619 : data_rom <= {16'd1943, 16'd32710};
                15'd620 : data_rom <= {16'd1946, 16'd32710};
                15'd621 : data_rom <= {16'd1949, 16'd32709};
                15'd622 : data_rom <= {16'd1952, 16'd32709};
                15'd623 : data_rom <= {16'd1956, 16'd32709};
                15'd624 : data_rom <= {16'd1959, 16'd32709};
                15'd625 : data_rom <= {16'd1962, 16'd32709};
                15'd626 : data_rom <= {16'd1965, 16'd32709};
                15'd627 : data_rom <= {16'd1968, 16'd32708};
                15'd628 : data_rom <= {16'd1971, 16'd32708};
                15'd629 : data_rom <= {16'd1974, 16'd32708};
                15'd630 : data_rom <= {16'd1977, 16'd32708};
                15'd631 : data_rom <= {16'd1981, 16'd32708};
                15'd632 : data_rom <= {16'd1984, 16'd32707};
                15'd633 : data_rom <= {16'd1987, 16'd32707};
                15'd634 : data_rom <= {16'd1990, 16'd32707};
                15'd635 : data_rom <= {16'd1993, 16'd32707};
                15'd636 : data_rom <= {16'd1996, 16'd32707};
                15'd637 : data_rom <= {16'd1999, 16'd32706};
                15'd638 : data_rom <= {16'd2003, 16'd32706};
                15'd639 : data_rom <= {16'd2006, 16'd32706};
                15'd640 : data_rom <= {16'd2009, 16'd32706};
                15'd641 : data_rom <= {16'd2012, 16'd32706};
                15'd642 : data_rom <= {16'd2015, 16'd32705};
                15'd643 : data_rom <= {16'd2018, 16'd32705};
                15'd644 : data_rom <= {16'd2021, 16'd32705};
                15'd645 : data_rom <= {16'd2025, 16'd32705};
                15'd646 : data_rom <= {16'd2028, 16'd32705};
                15'd647 : data_rom <= {16'd2031, 16'd32704};
                15'd648 : data_rom <= {16'd2034, 16'd32704};
                15'd649 : data_rom <= {16'd2037, 16'd32704};
                15'd650 : data_rom <= {16'd2040, 16'd32704};
                15'd651 : data_rom <= {16'd2043, 16'd32704};
                15'd652 : data_rom <= {16'd2046, 16'd32704};
                15'd653 : data_rom <= {16'd2050, 16'd32703};
                15'd654 : data_rom <= {16'd2053, 16'd32703};
                15'd655 : data_rom <= {16'd2056, 16'd32703};
                15'd656 : data_rom <= {16'd2059, 16'd32703};
                15'd657 : data_rom <= {16'd2062, 16'd32703};
                15'd658 : data_rom <= {16'd2065, 16'd32702};
                15'd659 : data_rom <= {16'd2068, 16'd32702};
                15'd660 : data_rom <= {16'd2072, 16'd32702};
                15'd661 : data_rom <= {16'd2075, 16'd32702};
                15'd662 : data_rom <= {16'd2078, 16'd32702};
                15'd663 : data_rom <= {16'd2081, 16'd32701};
                15'd664 : data_rom <= {16'd2084, 16'd32701};
                15'd665 : data_rom <= {16'd2087, 16'd32701};
                15'd666 : data_rom <= {16'd2090, 16'd32701};
                15'd667 : data_rom <= {16'd2094, 16'd32701};
                15'd668 : data_rom <= {16'd2097, 16'd32700};
                15'd669 : data_rom <= {16'd2100, 16'd32700};
                15'd670 : data_rom <= {16'd2103, 16'd32700};
                15'd671 : data_rom <= {16'd2106, 16'd32700};
                15'd672 : data_rom <= {16'd2109, 16'd32700};
                15'd673 : data_rom <= {16'd2112, 16'd32699};
                15'd674 : data_rom <= {16'd2115, 16'd32699};
                15'd675 : data_rom <= {16'd2119, 16'd32699};
                15'd676 : data_rom <= {16'd2122, 16'd32699};
                15'd677 : data_rom <= {16'd2125, 16'd32699};
                15'd678 : data_rom <= {16'd2128, 16'd32698};
                15'd679 : data_rom <= {16'd2131, 16'd32698};
                15'd680 : data_rom <= {16'd2134, 16'd32698};
                15'd681 : data_rom <= {16'd2137, 16'd32698};
                15'd682 : data_rom <= {16'd2141, 16'd32697};
                15'd683 : data_rom <= {16'd2144, 16'd32697};
                15'd684 : data_rom <= {16'd2147, 16'd32697};
                15'd685 : data_rom <= {16'd2150, 16'd32697};
                15'd686 : data_rom <= {16'd2153, 16'd32697};
                15'd687 : data_rom <= {16'd2156, 16'd32696};
                15'd688 : data_rom <= {16'd2159, 16'd32696};
                15'd689 : data_rom <= {16'd2162, 16'd32696};
                15'd690 : data_rom <= {16'd2166, 16'd32696};
                15'd691 : data_rom <= {16'd2169, 16'd32696};
                15'd692 : data_rom <= {16'd2172, 16'd32695};
                15'd693 : data_rom <= {16'd2175, 16'd32695};
                15'd694 : data_rom <= {16'd2178, 16'd32695};
                15'd695 : data_rom <= {16'd2181, 16'd32695};
                15'd696 : data_rom <= {16'd2184, 16'd32695};
                15'd697 : data_rom <= {16'd2188, 16'd32694};
                15'd698 : data_rom <= {16'd2191, 16'd32694};
                15'd699 : data_rom <= {16'd2194, 16'd32694};
                15'd700 : data_rom <= {16'd2197, 16'd32694};
                15'd701 : data_rom <= {16'd2200, 16'd32694};
                15'd702 : data_rom <= {16'd2203, 16'd32693};
                15'd703 : data_rom <= {16'd2206, 16'd32693};
                15'd704 : data_rom <= {16'd2210, 16'd32693};
                15'd705 : data_rom <= {16'd2213, 16'd32693};
                15'd706 : data_rom <= {16'd2216, 16'd32692};
                15'd707 : data_rom <= {16'd2219, 16'd32692};
                15'd708 : data_rom <= {16'd2222, 16'd32692};
                15'd709 : data_rom <= {16'd2225, 16'd32692};
                15'd710 : data_rom <= {16'd2228, 16'd32692};
                15'd711 : data_rom <= {16'd2231, 16'd32691};
                15'd712 : data_rom <= {16'd2235, 16'd32691};
                15'd713 : data_rom <= {16'd2238, 16'd32691};
                15'd714 : data_rom <= {16'd2241, 16'd32691};
                15'd715 : data_rom <= {16'd2244, 16'd32691};
                15'd716 : data_rom <= {16'd2247, 16'd32690};
                15'd717 : data_rom <= {16'd2250, 16'd32690};
                15'd718 : data_rom <= {16'd2253, 16'd32690};
                15'd719 : data_rom <= {16'd2257, 16'd32690};
                15'd720 : data_rom <= {16'd2260, 16'd32689};
                15'd721 : data_rom <= {16'd2263, 16'd32689};
                15'd722 : data_rom <= {16'd2266, 16'd32689};
                15'd723 : data_rom <= {16'd2269, 16'd32689};
                15'd724 : data_rom <= {16'd2272, 16'd32689};
                15'd725 : data_rom <= {16'd2275, 16'd32688};
                15'd726 : data_rom <= {16'd2278, 16'd32688};
                15'd727 : data_rom <= {16'd2282, 16'd32688};
                15'd728 : data_rom <= {16'd2285, 16'd32688};
                15'd729 : data_rom <= {16'd2288, 16'd32687};
                15'd730 : data_rom <= {16'd2291, 16'd32687};
                15'd731 : data_rom <= {16'd2294, 16'd32687};
                15'd732 : data_rom <= {16'd2297, 16'd32687};
                15'd733 : data_rom <= {16'd2300, 16'd32687};
                15'd734 : data_rom <= {16'd2304, 16'd32686};
                15'd735 : data_rom <= {16'd2307, 16'd32686};
                15'd736 : data_rom <= {16'd2310, 16'd32686};
                15'd737 : data_rom <= {16'd2313, 16'd32686};
                15'd738 : data_rom <= {16'd2316, 16'd32686};
                15'd739 : data_rom <= {16'd2319, 16'd32685};
                15'd740 : data_rom <= {16'd2322, 16'd32685};
                15'd741 : data_rom <= {16'd2325, 16'd32685};
                15'd742 : data_rom <= {16'd2329, 16'd32685};
                15'd743 : data_rom <= {16'd2332, 16'd32684};
                15'd744 : data_rom <= {16'd2335, 16'd32684};
                15'd745 : data_rom <= {16'd2338, 16'd32684};
                15'd746 : data_rom <= {16'd2341, 16'd32684};
                15'd747 : data_rom <= {16'd2344, 16'd32684};
                15'd748 : data_rom <= {16'd2347, 16'd32683};
                15'd749 : data_rom <= {16'd2351, 16'd32683};
                15'd750 : data_rom <= {16'd2354, 16'd32683};
                15'd751 : data_rom <= {16'd2357, 16'd32683};
                15'd752 : data_rom <= {16'd2360, 16'd32682};
                15'd753 : data_rom <= {16'd2363, 16'd32682};
                15'd754 : data_rom <= {16'd2366, 16'd32682};
                15'd755 : data_rom <= {16'd2369, 16'd32682};
                15'd756 : data_rom <= {16'd2372, 16'd32681};
                15'd757 : data_rom <= {16'd2376, 16'd32681};
                15'd758 : data_rom <= {16'd2379, 16'd32681};
                15'd759 : data_rom <= {16'd2382, 16'd32681};
                15'd760 : data_rom <= {16'd2385, 16'd32681};
                15'd761 : data_rom <= {16'd2388, 16'd32680};
                15'd762 : data_rom <= {16'd2391, 16'd32680};
                15'd763 : data_rom <= {16'd2394, 16'd32680};
                15'd764 : data_rom <= {16'd2398, 16'd32680};
                15'd765 : data_rom <= {16'd2401, 16'd32679};
                15'd766 : data_rom <= {16'd2404, 16'd32679};
                15'd767 : data_rom <= {16'd2407, 16'd32679};
                15'd768 : data_rom <= {16'd2410, 16'd32679};
                15'd769 : data_rom <= {16'd2413, 16'd32678};
                15'd770 : data_rom <= {16'd2416, 16'd32678};
                15'd771 : data_rom <= {16'd2419, 16'd32678};
                15'd772 : data_rom <= {16'd2423, 16'd32678};
                15'd773 : data_rom <= {16'd2426, 16'd32678};
                15'd774 : data_rom <= {16'd2429, 16'd32677};
                15'd775 : data_rom <= {16'd2432, 16'd32677};
                15'd776 : data_rom <= {16'd2435, 16'd32677};
                15'd777 : data_rom <= {16'd2438, 16'd32677};
                15'd778 : data_rom <= {16'd2441, 16'd32676};
                15'd779 : data_rom <= {16'd2445, 16'd32676};
                15'd780 : data_rom <= {16'd2448, 16'd32676};
                15'd781 : data_rom <= {16'd2451, 16'd32676};
                15'd782 : data_rom <= {16'd2454, 16'd32675};
                15'd783 : data_rom <= {16'd2457, 16'd32675};
                15'd784 : data_rom <= {16'd2460, 16'd32675};
                15'd785 : data_rom <= {16'd2463, 16'd32675};
                15'd786 : data_rom <= {16'd2466, 16'd32675};
                15'd787 : data_rom <= {16'd2470, 16'd32674};
                15'd788 : data_rom <= {16'd2473, 16'd32674};
                15'd789 : data_rom <= {16'd2476, 16'd32674};
                15'd790 : data_rom <= {16'd2479, 16'd32674};
                15'd791 : data_rom <= {16'd2482, 16'd32673};
                15'd792 : data_rom <= {16'd2485, 16'd32673};
                15'd793 : data_rom <= {16'd2488, 16'd32673};
                15'd794 : data_rom <= {16'd2492, 16'd32673};
                15'd795 : data_rom <= {16'd2495, 16'd32672};
                15'd796 : data_rom <= {16'd2498, 16'd32672};
                15'd797 : data_rom <= {16'd2501, 16'd32672};
                15'd798 : data_rom <= {16'd2504, 16'd32672};
                15'd799 : data_rom <= {16'd2507, 16'd32671};
                15'd800 : data_rom <= {16'd2510, 16'd32671};
                15'd801 : data_rom <= {16'd2513, 16'd32671};
                15'd802 : data_rom <= {16'd2517, 16'd32671};
                15'd803 : data_rom <= {16'd2520, 16'd32670};
                15'd804 : data_rom <= {16'd2523, 16'd32670};
                15'd805 : data_rom <= {16'd2526, 16'd32670};
                15'd806 : data_rom <= {16'd2529, 16'd32670};
                15'd807 : data_rom <= {16'd2532, 16'd32669};
                15'd808 : data_rom <= {16'd2535, 16'd32669};
                15'd809 : data_rom <= {16'd2538, 16'd32669};
                15'd810 : data_rom <= {16'd2542, 16'd32669};
                15'd811 : data_rom <= {16'd2545, 16'd32668};
                15'd812 : data_rom <= {16'd2548, 16'd32668};
                15'd813 : data_rom <= {16'd2551, 16'd32668};
                15'd814 : data_rom <= {16'd2554, 16'd32668};
                15'd815 : data_rom <= {16'd2557, 16'd32668};
                15'd816 : data_rom <= {16'd2560, 16'd32667};
                15'd817 : data_rom <= {16'd2564, 16'd32667};
                15'd818 : data_rom <= {16'd2567, 16'd32667};
                15'd819 : data_rom <= {16'd2570, 16'd32667};
                15'd820 : data_rom <= {16'd2573, 16'd32666};
                15'd821 : data_rom <= {16'd2576, 16'd32666};
                15'd822 : data_rom <= {16'd2579, 16'd32666};
                15'd823 : data_rom <= {16'd2582, 16'd32666};
                15'd824 : data_rom <= {16'd2585, 16'd32665};
                15'd825 : data_rom <= {16'd2589, 16'd32665};
                15'd826 : data_rom <= {16'd2592, 16'd32665};
                15'd827 : data_rom <= {16'd2595, 16'd32665};
                15'd828 : data_rom <= {16'd2598, 16'd32664};
                15'd829 : data_rom <= {16'd2601, 16'd32664};
                15'd830 : data_rom <= {16'd2604, 16'd32664};
                15'd831 : data_rom <= {16'd2607, 16'd32664};
                15'd832 : data_rom <= {16'd2611, 16'd32663};
                15'd833 : data_rom <= {16'd2614, 16'd32663};
                15'd834 : data_rom <= {16'd2617, 16'd32663};
                15'd835 : data_rom <= {16'd2620, 16'd32663};
                15'd836 : data_rom <= {16'd2623, 16'd32662};
                15'd837 : data_rom <= {16'd2626, 16'd32662};
                15'd838 : data_rom <= {16'd2629, 16'd32662};
                15'd839 : data_rom <= {16'd2632, 16'd32662};
                15'd840 : data_rom <= {16'd2636, 16'd32661};
                15'd841 : data_rom <= {16'd2639, 16'd32661};
                15'd842 : data_rom <= {16'd2642, 16'd32661};
                15'd843 : data_rom <= {16'd2645, 16'd32661};
                15'd844 : data_rom <= {16'd2648, 16'd32660};
                15'd845 : data_rom <= {16'd2651, 16'd32660};
                15'd846 : data_rom <= {16'd2654, 16'd32660};
                15'd847 : data_rom <= {16'd2658, 16'd32660};
                15'd848 : data_rom <= {16'd2661, 16'd32659};
                15'd849 : data_rom <= {16'd2664, 16'd32659};
                15'd850 : data_rom <= {16'd2667, 16'd32659};
                15'd851 : data_rom <= {16'd2670, 16'd32658};
                15'd852 : data_rom <= {16'd2673, 16'd32658};
                15'd853 : data_rom <= {16'd2676, 16'd32658};
                15'd854 : data_rom <= {16'd2679, 16'd32658};
                15'd855 : data_rom <= {16'd2683, 16'd32657};
                15'd856 : data_rom <= {16'd2686, 16'd32657};
                15'd857 : data_rom <= {16'd2689, 16'd32657};
                15'd858 : data_rom <= {16'd2692, 16'd32657};
                15'd859 : data_rom <= {16'd2695, 16'd32656};
                15'd860 : data_rom <= {16'd2698, 16'd32656};
                15'd861 : data_rom <= {16'd2701, 16'd32656};
                15'd862 : data_rom <= {16'd2704, 16'd32656};
                15'd863 : data_rom <= {16'd2708, 16'd32655};
                15'd864 : data_rom <= {16'd2711, 16'd32655};
                15'd865 : data_rom <= {16'd2714, 16'd32655};
                15'd866 : data_rom <= {16'd2717, 16'd32655};
                15'd867 : data_rom <= {16'd2720, 16'd32654};
                15'd868 : data_rom <= {16'd2723, 16'd32654};
                15'd869 : data_rom <= {16'd2726, 16'd32654};
                15'd870 : data_rom <= {16'd2730, 16'd32654};
                15'd871 : data_rom <= {16'd2733, 16'd32653};
                15'd872 : data_rom <= {16'd2736, 16'd32653};
                15'd873 : data_rom <= {16'd2739, 16'd32653};
                15'd874 : data_rom <= {16'd2742, 16'd32653};
                15'd875 : data_rom <= {16'd2745, 16'd32652};
                15'd876 : data_rom <= {16'd2748, 16'd32652};
                15'd877 : data_rom <= {16'd2751, 16'd32652};
                15'd878 : data_rom <= {16'd2755, 16'd32651};
                15'd879 : data_rom <= {16'd2758, 16'd32651};
                15'd880 : data_rom <= {16'd2761, 16'd32651};
                15'd881 : data_rom <= {16'd2764, 16'd32651};
                15'd882 : data_rom <= {16'd2767, 16'd32650};
                15'd883 : data_rom <= {16'd2770, 16'd32650};
                15'd884 : data_rom <= {16'd2773, 16'd32650};
                15'd885 : data_rom <= {16'd2776, 16'd32650};
                15'd886 : data_rom <= {16'd2780, 16'd32649};
                15'd887 : data_rom <= {16'd2783, 16'd32649};
                15'd888 : data_rom <= {16'd2786, 16'd32649};
                15'd889 : data_rom <= {16'd2789, 16'd32649};
                15'd890 : data_rom <= {16'd2792, 16'd32648};
                15'd891 : data_rom <= {16'd2795, 16'd32648};
                15'd892 : data_rom <= {16'd2798, 16'd32648};
                15'd893 : data_rom <= {16'd2802, 16'd32647};
                15'd894 : data_rom <= {16'd2805, 16'd32647};
                15'd895 : data_rom <= {16'd2808, 16'd32647};
                15'd896 : data_rom <= {16'd2811, 16'd32647};
                15'd897 : data_rom <= {16'd2814, 16'd32646};
                15'd898 : data_rom <= {16'd2817, 16'd32646};
                15'd899 : data_rom <= {16'd2820, 16'd32646};
                15'd900 : data_rom <= {16'd2823, 16'd32646};
                15'd901 : data_rom <= {16'd2827, 16'd32645};
                15'd902 : data_rom <= {16'd2830, 16'd32645};
                15'd903 : data_rom <= {16'd2833, 16'd32645};
                15'd904 : data_rom <= {16'd2836, 16'd32645};
                15'd905 : data_rom <= {16'd2839, 16'd32644};
                15'd906 : data_rom <= {16'd2842, 16'd32644};
                15'd907 : data_rom <= {16'd2845, 16'd32644};
                15'd908 : data_rom <= {16'd2848, 16'd32643};
                15'd909 : data_rom <= {16'd2852, 16'd32643};
                15'd910 : data_rom <= {16'd2855, 16'd32643};
                15'd911 : data_rom <= {16'd2858, 16'd32643};
                15'd912 : data_rom <= {16'd2861, 16'd32642};
                15'd913 : data_rom <= {16'd2864, 16'd32642};
                15'd914 : data_rom <= {16'd2867, 16'd32642};
                15'd915 : data_rom <= {16'd2870, 16'd32641};
                15'd916 : data_rom <= {16'd2873, 16'd32641};
                15'd917 : data_rom <= {16'd2877, 16'd32641};
                15'd918 : data_rom <= {16'd2880, 16'd32641};
                15'd919 : data_rom <= {16'd2883, 16'd32640};
                15'd920 : data_rom <= {16'd2886, 16'd32640};
                15'd921 : data_rom <= {16'd2889, 16'd32640};
                15'd922 : data_rom <= {16'd2892, 16'd32640};
                15'd923 : data_rom <= {16'd2895, 16'd32639};
                15'd924 : data_rom <= {16'd2899, 16'd32639};
                15'd925 : data_rom <= {16'd2902, 16'd32639};
                15'd926 : data_rom <= {16'd2905, 16'd32638};
                15'd927 : data_rom <= {16'd2908, 16'd32638};
                15'd928 : data_rom <= {16'd2911, 16'd32638};
                15'd929 : data_rom <= {16'd2914, 16'd32638};
                15'd930 : data_rom <= {16'd2917, 16'd32637};
                15'd931 : data_rom <= {16'd2920, 16'd32637};
                15'd932 : data_rom <= {16'd2924, 16'd32637};
                15'd933 : data_rom <= {16'd2927, 16'd32636};
                15'd934 : data_rom <= {16'd2930, 16'd32636};
                15'd935 : data_rom <= {16'd2933, 16'd32636};
                15'd936 : data_rom <= {16'd2936, 16'd32636};
                15'd937 : data_rom <= {16'd2939, 16'd32635};
                15'd938 : data_rom <= {16'd2942, 16'd32635};
                15'd939 : data_rom <= {16'd2945, 16'd32635};
                15'd940 : data_rom <= {16'd2949, 16'd32635};
                15'd941 : data_rom <= {16'd2952, 16'd32634};
                15'd942 : data_rom <= {16'd2955, 16'd32634};
                15'd943 : data_rom <= {16'd2958, 16'd32634};
                15'd944 : data_rom <= {16'd2961, 16'd32633};
                15'd945 : data_rom <= {16'd2964, 16'd32633};
                15'd946 : data_rom <= {16'd2967, 16'd32633};
                15'd947 : data_rom <= {16'd2970, 16'd32633};
                15'd948 : data_rom <= {16'd2974, 16'd32632};
                15'd949 : data_rom <= {16'd2977, 16'd32632};
                15'd950 : data_rom <= {16'd2980, 16'd32632};
                15'd951 : data_rom <= {16'd2983, 16'd32631};
                15'd952 : data_rom <= {16'd2986, 16'd32631};
                15'd953 : data_rom <= {16'd2989, 16'd32631};
                15'd954 : data_rom <= {16'd2992, 16'd32631};
                15'd955 : data_rom <= {16'd2996, 16'd32630};
                15'd956 : data_rom <= {16'd2999, 16'd32630};
                15'd957 : data_rom <= {16'd3002, 16'd32630};
                15'd958 : data_rom <= {16'd3005, 16'd32629};
                15'd959 : data_rom <= {16'd3008, 16'd32629};
                15'd960 : data_rom <= {16'd3011, 16'd32629};
                15'd961 : data_rom <= {16'd3014, 16'd32629};
                15'd962 : data_rom <= {16'd3017, 16'd32628};
                15'd963 : data_rom <= {16'd3021, 16'd32628};
                15'd964 : data_rom <= {16'd3024, 16'd32628};
                15'd965 : data_rom <= {16'd3027, 16'd32627};
                15'd966 : data_rom <= {16'd3030, 16'd32627};
                15'd967 : data_rom <= {16'd3033, 16'd32627};
                15'd968 : data_rom <= {16'd3036, 16'd32626};
                15'd969 : data_rom <= {16'd3039, 16'd32626};
                15'd970 : data_rom <= {16'd3042, 16'd32626};
                15'd971 : data_rom <= {16'd3046, 16'd32626};
                15'd972 : data_rom <= {16'd3049, 16'd32625};
                15'd973 : data_rom <= {16'd3052, 16'd32625};
                15'd974 : data_rom <= {16'd3055, 16'd32625};
                15'd975 : data_rom <= {16'd3058, 16'd32624};
                15'd976 : data_rom <= {16'd3061, 16'd32624};
                15'd977 : data_rom <= {16'd3064, 16'd32624};
                15'd978 : data_rom <= {16'd3067, 16'd32624};
                15'd979 : data_rom <= {16'd3071, 16'd32623};
                15'd980 : data_rom <= {16'd3074, 16'd32623};
                15'd981 : data_rom <= {16'd3077, 16'd32623};
                15'd982 : data_rom <= {16'd3080, 16'd32622};
                15'd983 : data_rom <= {16'd3083, 16'd32622};
                15'd984 : data_rom <= {16'd3086, 16'd32622};
                15'd985 : data_rom <= {16'd3089, 16'd32621};
                15'd986 : data_rom <= {16'd3092, 16'd32621};
                15'd987 : data_rom <= {16'd3096, 16'd32621};
                15'd988 : data_rom <= {16'd3099, 16'd32621};
                15'd989 : data_rom <= {16'd3102, 16'd32620};
                15'd990 : data_rom <= {16'd3105, 16'd32620};
                15'd991 : data_rom <= {16'd3108, 16'd32620};
                15'd992 : data_rom <= {16'd3111, 16'd32619};
                15'd993 : data_rom <= {16'd3114, 16'd32619};
                15'd994 : data_rom <= {16'd3118, 16'd32619};
                15'd995 : data_rom <= {16'd3121, 16'd32619};
                15'd996 : data_rom <= {16'd3124, 16'd32618};
                15'd997 : data_rom <= {16'd3127, 16'd32618};
                15'd998 : data_rom <= {16'd3130, 16'd32618};
                15'd999 : data_rom <= {16'd3133, 16'd32617};
                15'd1000 : data_rom <= {16'd3136, 16'd32617};
                15'd1001 : data_rom <= {16'd3139, 16'd32617};
                15'd1002 : data_rom <= {16'd3143, 16'd32616};
                15'd1003 : data_rom <= {16'd3146, 16'd32616};
                15'd1004 : data_rom <= {16'd3149, 16'd32616};
                15'd1005 : data_rom <= {16'd3152, 16'd32616};
                15'd1006 : data_rom <= {16'd3155, 16'd32615};
                15'd1007 : data_rom <= {16'd3158, 16'd32615};
                15'd1008 : data_rom <= {16'd3161, 16'd32615};
                15'd1009 : data_rom <= {16'd3164, 16'd32614};
                15'd1010 : data_rom <= {16'd3168, 16'd32614};
                15'd1011 : data_rom <= {16'd3171, 16'd32614};
                15'd1012 : data_rom <= {16'd3174, 16'd32613};
                15'd1013 : data_rom <= {16'd3177, 16'd32613};
                15'd1014 : data_rom <= {16'd3180, 16'd32613};
                15'd1015 : data_rom <= {16'd3183, 16'd32612};
                15'd1016 : data_rom <= {16'd3186, 16'd32612};
                15'd1017 : data_rom <= {16'd3189, 16'd32612};
                15'd1018 : data_rom <= {16'd3193, 16'd32612};
                15'd1019 : data_rom <= {16'd3196, 16'd32611};
                15'd1020 : data_rom <= {16'd3199, 16'd32611};
                15'd1021 : data_rom <= {16'd3202, 16'd32611};
                15'd1022 : data_rom <= {16'd3205, 16'd32610};
                15'd1023 : data_rom <= {16'd3208, 16'd32610};
                15'd1024 : data_rom <= {16'd3211, 16'd32610};
                15'd1025 : data_rom <= {16'd3214, 16'd32609};
                15'd1026 : data_rom <= {16'd3218, 16'd32609};
                15'd1027 : data_rom <= {16'd3221, 16'd32609};
                15'd1028 : data_rom <= {16'd3224, 16'd32608};
                15'd1029 : data_rom <= {16'd3227, 16'd32608};
                15'd1030 : data_rom <= {16'd3230, 16'd32608};
                15'd1031 : data_rom <= {16'd3233, 16'd32608};
                15'd1032 : data_rom <= {16'd3236, 16'd32607};
                15'd1033 : data_rom <= {16'd3239, 16'd32607};
                15'd1034 : data_rom <= {16'd3243, 16'd32607};
                15'd1035 : data_rom <= {16'd3246, 16'd32606};
                15'd1036 : data_rom <= {16'd3249, 16'd32606};
                15'd1037 : data_rom <= {16'd3252, 16'd32606};
                15'd1038 : data_rom <= {16'd3255, 16'd32605};
                15'd1039 : data_rom <= {16'd3258, 16'd32605};
                15'd1040 : data_rom <= {16'd3261, 16'd32605};
                15'd1041 : data_rom <= {16'd3264, 16'd32604};
                15'd1042 : data_rom <= {16'd3268, 16'd32604};
                15'd1043 : data_rom <= {16'd3271, 16'd32604};
                15'd1044 : data_rom <= {16'd3274, 16'd32603};
                15'd1045 : data_rom <= {16'd3277, 16'd32603};
                15'd1046 : data_rom <= {16'd3280, 16'd32603};
                15'd1047 : data_rom <= {16'd3283, 16'd32603};
                15'd1048 : data_rom <= {16'd3286, 16'd32602};
                15'd1049 : data_rom <= {16'd3289, 16'd32602};
                15'd1050 : data_rom <= {16'd3293, 16'd32602};
                15'd1051 : data_rom <= {16'd3296, 16'd32601};
                15'd1052 : data_rom <= {16'd3299, 16'd32601};
                15'd1053 : data_rom <= {16'd3302, 16'd32601};
                15'd1054 : data_rom <= {16'd3305, 16'd32600};
                15'd1055 : data_rom <= {16'd3308, 16'd32600};
                15'd1056 : data_rom <= {16'd3311, 16'd32600};
                15'd1057 : data_rom <= {16'd3314, 16'd32599};
                15'd1058 : data_rom <= {16'd3318, 16'd32599};
                15'd1059 : data_rom <= {16'd3321, 16'd32599};
                15'd1060 : data_rom <= {16'd3324, 16'd32598};
                15'd1061 : data_rom <= {16'd3327, 16'd32598};
                15'd1062 : data_rom <= {16'd3330, 16'd32598};
                15'd1063 : data_rom <= {16'd3333, 16'd32597};
                15'd1064 : data_rom <= {16'd3336, 16'd32597};
                15'd1065 : data_rom <= {16'd3339, 16'd32597};
                15'd1066 : data_rom <= {16'd3343, 16'd32597};
                15'd1067 : data_rom <= {16'd3346, 16'd32596};
                15'd1068 : data_rom <= {16'd3349, 16'd32596};
                15'd1069 : data_rom <= {16'd3352, 16'd32596};
                15'd1070 : data_rom <= {16'd3355, 16'd32595};
                15'd1071 : data_rom <= {16'd3358, 16'd32595};
                15'd1072 : data_rom <= {16'd3361, 16'd32595};
                15'd1073 : data_rom <= {16'd3364, 16'd32594};
                15'd1074 : data_rom <= {16'd3368, 16'd32594};
                15'd1075 : data_rom <= {16'd3371, 16'd32594};
                15'd1076 : data_rom <= {16'd3374, 16'd32593};
                15'd1077 : data_rom <= {16'd3377, 16'd32593};
                15'd1078 : data_rom <= {16'd3380, 16'd32593};
                15'd1079 : data_rom <= {16'd3383, 16'd32592};
                15'd1080 : data_rom <= {16'd3386, 16'd32592};
                15'd1081 : data_rom <= {16'd3389, 16'd32592};
                15'd1082 : data_rom <= {16'd3393, 16'd32591};
                15'd1083 : data_rom <= {16'd3396, 16'd32591};
                15'd1084 : data_rom <= {16'd3399, 16'd32591};
                15'd1085 : data_rom <= {16'd3402, 16'd32590};
                15'd1086 : data_rom <= {16'd3405, 16'd32590};
                15'd1087 : data_rom <= {16'd3408, 16'd32590};
                15'd1088 : data_rom <= {16'd3411, 16'd32589};
                15'd1089 : data_rom <= {16'd3414, 16'd32589};
                15'd1090 : data_rom <= {16'd3418, 16'd32589};
                15'd1091 : data_rom <= {16'd3421, 16'd32588};
                15'd1092 : data_rom <= {16'd3424, 16'd32588};
                15'd1093 : data_rom <= {16'd3427, 16'd32588};
                15'd1094 : data_rom <= {16'd3430, 16'd32587};
                15'd1095 : data_rom <= {16'd3433, 16'd32587};
                15'd1096 : data_rom <= {16'd3436, 16'd32587};
                15'd1097 : data_rom <= {16'd3439, 16'd32586};
                15'd1098 : data_rom <= {16'd3443, 16'd32586};
                15'd1099 : data_rom <= {16'd3446, 16'd32586};
                15'd1100 : data_rom <= {16'd3449, 16'd32585};
                15'd1101 : data_rom <= {16'd3452, 16'd32585};
                15'd1102 : data_rom <= {16'd3455, 16'd32585};
                15'd1103 : data_rom <= {16'd3458, 16'd32584};
                15'd1104 : data_rom <= {16'd3461, 16'd32584};
                15'd1105 : data_rom <= {16'd3464, 16'd32584};
                15'd1106 : data_rom <= {16'd3468, 16'd32583};
                15'd1107 : data_rom <= {16'd3471, 16'd32583};
                15'd1108 : data_rom <= {16'd3474, 16'd32583};
                15'd1109 : data_rom <= {16'd3477, 16'd32582};
                15'd1110 : data_rom <= {16'd3480, 16'd32582};
                15'd1111 : data_rom <= {16'd3483, 16'd32582};
                15'd1112 : data_rom <= {16'd3486, 16'd32581};
                15'd1113 : data_rom <= {16'd3489, 16'd32581};
                15'd1114 : data_rom <= {16'd3493, 16'd32581};
                15'd1115 : data_rom <= {16'd3496, 16'd32580};
                15'd1116 : data_rom <= {16'd3499, 16'd32580};
                15'd1117 : data_rom <= {16'd3502, 16'd32580};
                15'd1118 : data_rom <= {16'd3505, 16'd32579};
                15'd1119 : data_rom <= {16'd3508, 16'd32579};
                15'd1120 : data_rom <= {16'd3511, 16'd32579};
                15'd1121 : data_rom <= {16'd3514, 16'd32578};
                15'd1122 : data_rom <= {16'd3518, 16'd32578};
                15'd1123 : data_rom <= {16'd3521, 16'd32578};
                15'd1124 : data_rom <= {16'd3524, 16'd32577};
                15'd1125 : data_rom <= {16'd3527, 16'd32577};
                15'd1126 : data_rom <= {16'd3530, 16'd32577};
                15'd1127 : data_rom <= {16'd3533, 16'd32576};
                15'd1128 : data_rom <= {16'd3536, 16'd32576};
                15'd1129 : data_rom <= {16'd3539, 16'd32576};
                15'd1130 : data_rom <= {16'd3543, 16'd32575};
                15'd1131 : data_rom <= {16'd3546, 16'd32575};
                15'd1132 : data_rom <= {16'd3549, 16'd32575};
                15'd1133 : data_rom <= {16'd3552, 16'd32574};
                15'd1134 : data_rom <= {16'd3555, 16'd32574};
                15'd1135 : data_rom <= {16'd3558, 16'd32574};
                15'd1136 : data_rom <= {16'd3561, 16'd32573};
                15'd1137 : data_rom <= {16'd3564, 16'd32573};
                15'd1138 : data_rom <= {16'd3568, 16'd32573};
                15'd1139 : data_rom <= {16'd3571, 16'd32572};
                15'd1140 : data_rom <= {16'd3574, 16'd32572};
                15'd1141 : data_rom <= {16'd3577, 16'd32572};
                15'd1142 : data_rom <= {16'd3580, 16'd32571};
                15'd1143 : data_rom <= {16'd3583, 16'd32571};
                15'd1144 : data_rom <= {16'd3586, 16'd32571};
                15'd1145 : data_rom <= {16'd3589, 16'd32570};
                15'd1146 : data_rom <= {16'd3593, 16'd32570};
                15'd1147 : data_rom <= {16'd3596, 16'd32570};
                15'd1148 : data_rom <= {16'd3599, 16'd32569};
                15'd1149 : data_rom <= {16'd3602, 16'd32569};
                15'd1150 : data_rom <= {16'd3605, 16'd32569};
                15'd1151 : data_rom <= {16'd3608, 16'd32568};
                15'd1152 : data_rom <= {16'd3611, 16'd32568};
                15'd1153 : data_rom <= {16'd3614, 16'd32567};
                15'd1154 : data_rom <= {16'd3618, 16'd32567};
                15'd1155 : data_rom <= {16'd3621, 16'd32567};
                15'd1156 : data_rom <= {16'd3624, 16'd32566};
                15'd1157 : data_rom <= {16'd3627, 16'd32566};
                15'd1158 : data_rom <= {16'd3630, 16'd32566};
                15'd1159 : data_rom <= {16'd3633, 16'd32565};
                15'd1160 : data_rom <= {16'd3636, 16'd32565};
                15'd1161 : data_rom <= {16'd3639, 16'd32565};
                15'd1162 : data_rom <= {16'd3642, 16'd32564};
                15'd1163 : data_rom <= {16'd3646, 16'd32564};
                15'd1164 : data_rom <= {16'd3649, 16'd32564};
                15'd1165 : data_rom <= {16'd3652, 16'd32563};
                15'd1166 : data_rom <= {16'd3655, 16'd32563};
                15'd1167 : data_rom <= {16'd3658, 16'd32563};
                15'd1168 : data_rom <= {16'd3661, 16'd32562};
                15'd1169 : data_rom <= {16'd3664, 16'd32562};
                15'd1170 : data_rom <= {16'd3667, 16'd32562};
                15'd1171 : data_rom <= {16'd3671, 16'd32561};
                15'd1172 : data_rom <= {16'd3674, 16'd32561};
                15'd1173 : data_rom <= {16'd3677, 16'd32561};
                15'd1174 : data_rom <= {16'd3680, 16'd32560};
                15'd1175 : data_rom <= {16'd3683, 16'd32560};
                15'd1176 : data_rom <= {16'd3686, 16'd32559};
                15'd1177 : data_rom <= {16'd3689, 16'd32559};
                15'd1178 : data_rom <= {16'd3692, 16'd32559};
                15'd1179 : data_rom <= {16'd3696, 16'd32558};
                15'd1180 : data_rom <= {16'd3699, 16'd32558};
                15'd1181 : data_rom <= {16'd3702, 16'd32558};
                15'd1182 : data_rom <= {16'd3705, 16'd32557};
                15'd1183 : data_rom <= {16'd3708, 16'd32557};
                15'd1184 : data_rom <= {16'd3711, 16'd32557};
                15'd1185 : data_rom <= {16'd3714, 16'd32556};
                15'd1186 : data_rom <= {16'd3717, 16'd32556};
                15'd1187 : data_rom <= {16'd3721, 16'd32556};
                15'd1188 : data_rom <= {16'd3724, 16'd32555};
                15'd1189 : data_rom <= {16'd3727, 16'd32555};
                15'd1190 : data_rom <= {16'd3730, 16'd32554};
                15'd1191 : data_rom <= {16'd3733, 16'd32554};
                15'd1192 : data_rom <= {16'd3736, 16'd32554};
                15'd1193 : data_rom <= {16'd3739, 16'd32553};
                15'd1194 : data_rom <= {16'd3742, 16'd32553};
                15'd1195 : data_rom <= {16'd3745, 16'd32553};
                15'd1196 : data_rom <= {16'd3749, 16'd32552};
                15'd1197 : data_rom <= {16'd3752, 16'd32552};
                15'd1198 : data_rom <= {16'd3755, 16'd32552};
                15'd1199 : data_rom <= {16'd3758, 16'd32551};
                15'd1200 : data_rom <= {16'd3761, 16'd32551};
                15'd1201 : data_rom <= {16'd3764, 16'd32551};
                15'd1202 : data_rom <= {16'd3767, 16'd32550};
                15'd1203 : data_rom <= {16'd3770, 16'd32550};
                15'd1204 : data_rom <= {16'd3774, 16'd32549};
                15'd1205 : data_rom <= {16'd3777, 16'd32549};
                15'd1206 : data_rom <= {16'd3780, 16'd32549};
                15'd1207 : data_rom <= {16'd3783, 16'd32548};
                15'd1208 : data_rom <= {16'd3786, 16'd32548};
                15'd1209 : data_rom <= {16'd3789, 16'd32548};
                15'd1210 : data_rom <= {16'd3792, 16'd32547};
                15'd1211 : data_rom <= {16'd3795, 16'd32547};
                15'd1212 : data_rom <= {16'd3799, 16'd32547};
                15'd1213 : data_rom <= {16'd3802, 16'd32546};
                15'd1214 : data_rom <= {16'd3805, 16'd32546};
                15'd1215 : data_rom <= {16'd3808, 16'd32545};
                15'd1216 : data_rom <= {16'd3811, 16'd32545};
                15'd1217 : data_rom <= {16'd3814, 16'd32545};
                15'd1218 : data_rom <= {16'd3817, 16'd32544};
                15'd1219 : data_rom <= {16'd3820, 16'd32544};
                15'd1220 : data_rom <= {16'd3824, 16'd32544};
                15'd1221 : data_rom <= {16'd3827, 16'd32543};
                15'd1222 : data_rom <= {16'd3830, 16'd32543};
                15'd1223 : data_rom <= {16'd3833, 16'd32543};
                15'd1224 : data_rom <= {16'd3836, 16'd32542};
                15'd1225 : data_rom <= {16'd3839, 16'd32542};
                15'd1226 : data_rom <= {16'd3842, 16'd32541};
                15'd1227 : data_rom <= {16'd3845, 16'd32541};
                15'd1228 : data_rom <= {16'd3848, 16'd32541};
                15'd1229 : data_rom <= {16'd3852, 16'd32540};
                15'd1230 : data_rom <= {16'd3855, 16'd32540};
                15'd1231 : data_rom <= {16'd3858, 16'd32540};
                15'd1232 : data_rom <= {16'd3861, 16'd32539};
                15'd1233 : data_rom <= {16'd3864, 16'd32539};
                15'd1234 : data_rom <= {16'd3867, 16'd32538};
                15'd1235 : data_rom <= {16'd3870, 16'd32538};
                15'd1236 : data_rom <= {16'd3873, 16'd32538};
                15'd1237 : data_rom <= {16'd3877, 16'd32537};
                15'd1238 : data_rom <= {16'd3880, 16'd32537};
                15'd1239 : data_rom <= {16'd3883, 16'd32537};
                15'd1240 : data_rom <= {16'd3886, 16'd32536};
                15'd1241 : data_rom <= {16'd3889, 16'd32536};
                15'd1242 : data_rom <= {16'd3892, 16'd32535};
                15'd1243 : data_rom <= {16'd3895, 16'd32535};
                15'd1244 : data_rom <= {16'd3898, 16'd32535};
                15'd1245 : data_rom <= {16'd3901, 16'd32534};
                15'd1246 : data_rom <= {16'd3905, 16'd32534};
                15'd1247 : data_rom <= {16'd3908, 16'd32534};
                15'd1248 : data_rom <= {16'd3911, 16'd32533};
                15'd1249 : data_rom <= {16'd3914, 16'd32533};
                15'd1250 : data_rom <= {16'd3917, 16'd32532};
                15'd1251 : data_rom <= {16'd3920, 16'd32532};
                15'd1252 : data_rom <= {16'd3923, 16'd32532};
                15'd1253 : data_rom <= {16'd3926, 16'd32531};
                15'd1254 : data_rom <= {16'd3930, 16'd32531};
                15'd1255 : data_rom <= {16'd3933, 16'd32531};
                15'd1256 : data_rom <= {16'd3936, 16'd32530};
                15'd1257 : data_rom <= {16'd3939, 16'd32530};
                15'd1258 : data_rom <= {16'd3942, 16'd32529};
                15'd1259 : data_rom <= {16'd3945, 16'd32529};
                15'd1260 : data_rom <= {16'd3948, 16'd32529};
                15'd1261 : data_rom <= {16'd3951, 16'd32528};
                15'd1262 : data_rom <= {16'd3955, 16'd32528};
                15'd1263 : data_rom <= {16'd3958, 16'd32528};
                15'd1264 : data_rom <= {16'd3961, 16'd32527};
                15'd1265 : data_rom <= {16'd3964, 16'd32527};
                15'd1266 : data_rom <= {16'd3967, 16'd32526};
                15'd1267 : data_rom <= {16'd3970, 16'd32526};
                15'd1268 : data_rom <= {16'd3973, 16'd32526};
                15'd1269 : data_rom <= {16'd3976, 16'd32525};
                15'd1270 : data_rom <= {16'd3979, 16'd32525};
                15'd1271 : data_rom <= {16'd3983, 16'd32525};
                15'd1272 : data_rom <= {16'd3986, 16'd32524};
                15'd1273 : data_rom <= {16'd3989, 16'd32524};
                15'd1274 : data_rom <= {16'd3992, 16'd32523};
                15'd1275 : data_rom <= {16'd3995, 16'd32523};
                15'd1276 : data_rom <= {16'd3998, 16'd32523};
                15'd1277 : data_rom <= {16'd4001, 16'd32522};
                15'd1278 : data_rom <= {16'd4004, 16'd32522};
                15'd1279 : data_rom <= {16'd4008, 16'd32521};
                15'd1280 : data_rom <= {16'd4011, 16'd32521};
                15'd1281 : data_rom <= {16'd4014, 16'd32521};
                15'd1282 : data_rom <= {16'd4017, 16'd32520};
                15'd1283 : data_rom <= {16'd4020, 16'd32520};
                15'd1284 : data_rom <= {16'd4023, 16'd32520};
                15'd1285 : data_rom <= {16'd4026, 16'd32519};
                15'd1286 : data_rom <= {16'd4029, 16'd32519};
                15'd1287 : data_rom <= {16'd4032, 16'd32518};
                15'd1288 : data_rom <= {16'd4036, 16'd32518};
                15'd1289 : data_rom <= {16'd4039, 16'd32518};
                15'd1290 : data_rom <= {16'd4042, 16'd32517};
                15'd1291 : data_rom <= {16'd4045, 16'd32517};
                15'd1292 : data_rom <= {16'd4048, 16'd32516};
                15'd1293 : data_rom <= {16'd4051, 16'd32516};
                15'd1294 : data_rom <= {16'd4054, 16'd32516};
                15'd1295 : data_rom <= {16'd4057, 16'd32515};
                15'd1296 : data_rom <= {16'd4061, 16'd32515};
                15'd1297 : data_rom <= {16'd4064, 16'd32514};
                15'd1298 : data_rom <= {16'd4067, 16'd32514};
                15'd1299 : data_rom <= {16'd4070, 16'd32514};
                15'd1300 : data_rom <= {16'd4073, 16'd32513};
                15'd1301 : data_rom <= {16'd4076, 16'd32513};
                15'd1302 : data_rom <= {16'd4079, 16'd32513};
                15'd1303 : data_rom <= {16'd4082, 16'd32512};
                15'd1304 : data_rom <= {16'd4085, 16'd32512};
                15'd1305 : data_rom <= {16'd4089, 16'd32511};
                15'd1306 : data_rom <= {16'd4092, 16'd32511};
                15'd1307 : data_rom <= {16'd4095, 16'd32511};
                15'd1308 : data_rom <= {16'd4098, 16'd32510};
                15'd1309 : data_rom <= {16'd4101, 16'd32510};
                15'd1310 : data_rom <= {16'd4104, 16'd32509};
                15'd1311 : data_rom <= {16'd4107, 16'd32509};
                15'd1312 : data_rom <= {16'd4110, 16'd32509};
                15'd1313 : data_rom <= {16'd4114, 16'd32508};
                15'd1314 : data_rom <= {16'd4117, 16'd32508};
                15'd1315 : data_rom <= {16'd4120, 16'd32507};
                15'd1316 : data_rom <= {16'd4123, 16'd32507};
                15'd1317 : data_rom <= {16'd4126, 16'd32507};
                15'd1318 : data_rom <= {16'd4129, 16'd32506};
                15'd1319 : data_rom <= {16'd4132, 16'd32506};
                15'd1320 : data_rom <= {16'd4135, 16'd32505};
                15'd1321 : data_rom <= {16'd4138, 16'd32505};
                15'd1322 : data_rom <= {16'd4142, 16'd32505};
                15'd1323 : data_rom <= {16'd4145, 16'd32504};
                15'd1324 : data_rom <= {16'd4148, 16'd32504};
                15'd1325 : data_rom <= {16'd4151, 16'd32503};
                15'd1326 : data_rom <= {16'd4154, 16'd32503};
                15'd1327 : data_rom <= {16'd4157, 16'd32503};
                15'd1328 : data_rom <= {16'd4160, 16'd32502};
                15'd1329 : data_rom <= {16'd4163, 16'd32502};
                15'd1330 : data_rom <= {16'd4167, 16'd32501};
                15'd1331 : data_rom <= {16'd4170, 16'd32501};
                15'd1332 : data_rom <= {16'd4173, 16'd32501};
                15'd1333 : data_rom <= {16'd4176, 16'd32500};
                15'd1334 : data_rom <= {16'd4179, 16'd32500};
                15'd1335 : data_rom <= {16'd4182, 16'd32499};
                15'd1336 : data_rom <= {16'd4185, 16'd32499};
                15'd1337 : data_rom <= {16'd4188, 16'd32499};
                15'd1338 : data_rom <= {16'd4191, 16'd32498};
                15'd1339 : data_rom <= {16'd4195, 16'd32498};
                15'd1340 : data_rom <= {16'd4198, 16'd32497};
                15'd1341 : data_rom <= {16'd4201, 16'd32497};
                15'd1342 : data_rom <= {16'd4204, 16'd32497};
                15'd1343 : data_rom <= {16'd4207, 16'd32496};
                15'd1344 : data_rom <= {16'd4210, 16'd32496};
                15'd1345 : data_rom <= {16'd4213, 16'd32495};
                15'd1346 : data_rom <= {16'd4216, 16'd32495};
                15'd1347 : data_rom <= {16'd4219, 16'd32495};
                15'd1348 : data_rom <= {16'd4223, 16'd32494};
                15'd1349 : data_rom <= {16'd4226, 16'd32494};
                15'd1350 : data_rom <= {16'd4229, 16'd32493};
                15'd1351 : data_rom <= {16'd4232, 16'd32493};
                15'd1352 : data_rom <= {16'd4235, 16'd32493};
                15'd1353 : data_rom <= {16'd4238, 16'd32492};
                15'd1354 : data_rom <= {16'd4241, 16'd32492};
                15'd1355 : data_rom <= {16'd4244, 16'd32491};
                15'd1356 : data_rom <= {16'd4248, 16'd32491};
                15'd1357 : data_rom <= {16'd4251, 16'd32491};
                15'd1358 : data_rom <= {16'd4254, 16'd32490};
                15'd1359 : data_rom <= {16'd4257, 16'd32490};
                15'd1360 : data_rom <= {16'd4260, 16'd32489};
                15'd1361 : data_rom <= {16'd4263, 16'd32489};
                15'd1362 : data_rom <= {16'd4266, 16'd32489};
                15'd1363 : data_rom <= {16'd4269, 16'd32488};
                15'd1364 : data_rom <= {16'd4272, 16'd32488};
                15'd1365 : data_rom <= {16'd4276, 16'd32487};
                15'd1366 : data_rom <= {16'd4279, 16'd32487};
                15'd1367 : data_rom <= {16'd4282, 16'd32486};
                15'd1368 : data_rom <= {16'd4285, 16'd32486};
                15'd1369 : data_rom <= {16'd4288, 16'd32486};
                15'd1370 : data_rom <= {16'd4291, 16'd32485};
                15'd1371 : data_rom <= {16'd4294, 16'd32485};
                15'd1372 : data_rom <= {16'd4297, 16'd32484};
                15'd1373 : data_rom <= {16'd4300, 16'd32484};
                15'd1374 : data_rom <= {16'd4304, 16'd32484};
                15'd1375 : data_rom <= {16'd4307, 16'd32483};
                15'd1376 : data_rom <= {16'd4310, 16'd32483};
                15'd1377 : data_rom <= {16'd4313, 16'd32482};
                15'd1378 : data_rom <= {16'd4316, 16'd32482};
                15'd1379 : data_rom <= {16'd4319, 16'd32482};
                15'd1380 : data_rom <= {16'd4322, 16'd32481};
                15'd1381 : data_rom <= {16'd4325, 16'd32481};
                15'd1382 : data_rom <= {16'd4328, 16'd32480};
                15'd1383 : data_rom <= {16'd4332, 16'd32480};
                15'd1384 : data_rom <= {16'd4335, 16'd32479};
                15'd1385 : data_rom <= {16'd4338, 16'd32479};
                15'd1386 : data_rom <= {16'd4341, 16'd32479};
                15'd1387 : data_rom <= {16'd4344, 16'd32478};
                15'd1388 : data_rom <= {16'd4347, 16'd32478};
                15'd1389 : data_rom <= {16'd4350, 16'd32477};
                15'd1390 : data_rom <= {16'd4353, 16'd32477};
                15'd1391 : data_rom <= {16'd4357, 16'd32477};
                15'd1392 : data_rom <= {16'd4360, 16'd32476};
                15'd1393 : data_rom <= {16'd4363, 16'd32476};
                15'd1394 : data_rom <= {16'd4366, 16'd32475};
                15'd1395 : data_rom <= {16'd4369, 16'd32475};
                15'd1396 : data_rom <= {16'd4372, 16'd32474};
                15'd1397 : data_rom <= {16'd4375, 16'd32474};
                15'd1398 : data_rom <= {16'd4378, 16'd32474};
                15'd1399 : data_rom <= {16'd4381, 16'd32473};
                15'd1400 : data_rom <= {16'd4385, 16'd32473};
                15'd1401 : data_rom <= {16'd4388, 16'd32472};
                15'd1402 : data_rom <= {16'd4391, 16'd32472};
                15'd1403 : data_rom <= {16'd4394, 16'd32472};
                15'd1404 : data_rom <= {16'd4397, 16'd32471};
                15'd1405 : data_rom <= {16'd4400, 16'd32471};
                15'd1406 : data_rom <= {16'd4403, 16'd32470};
                15'd1407 : data_rom <= {16'd4406, 16'd32470};
                15'd1408 : data_rom <= {16'd4409, 16'd32469};
                15'd1409 : data_rom <= {16'd4413, 16'd32469};
                15'd1410 : data_rom <= {16'd4416, 16'd32469};
                15'd1411 : data_rom <= {16'd4419, 16'd32468};
                15'd1412 : data_rom <= {16'd4422, 16'd32468};
                15'd1413 : data_rom <= {16'd4425, 16'd32467};
                15'd1414 : data_rom <= {16'd4428, 16'd32467};
                15'd1415 : data_rom <= {16'd4431, 16'd32466};
                15'd1416 : data_rom <= {16'd4434, 16'd32466};
                15'd1417 : data_rom <= {16'd4437, 16'd32466};
                15'd1418 : data_rom <= {16'd4441, 16'd32465};
                15'd1419 : data_rom <= {16'd4444, 16'd32465};
                15'd1420 : data_rom <= {16'd4447, 16'd32464};
                15'd1421 : data_rom <= {16'd4450, 16'd32464};
                15'd1422 : data_rom <= {16'd4453, 16'd32463};
                15'd1423 : data_rom <= {16'd4456, 16'd32463};
                15'd1424 : data_rom <= {16'd4459, 16'd32463};
                15'd1425 : data_rom <= {16'd4462, 16'd32462};
                15'd1426 : data_rom <= {16'd4465, 16'd32462};
                15'd1427 : data_rom <= {16'd4469, 16'd32461};
                15'd1428 : data_rom <= {16'd4472, 16'd32461};
                15'd1429 : data_rom <= {16'd4475, 16'd32460};
                15'd1430 : data_rom <= {16'd4478, 16'd32460};
                15'd1431 : data_rom <= {16'd4481, 16'd32460};
                15'd1432 : data_rom <= {16'd4484, 16'd32459};
                15'd1433 : data_rom <= {16'd4487, 16'd32459};
                15'd1434 : data_rom <= {16'd4490, 16'd32458};
                15'd1435 : data_rom <= {16'd4493, 16'd32458};
                15'd1436 : data_rom <= {16'd4497, 16'd32457};
                15'd1437 : data_rom <= {16'd4500, 16'd32457};
                15'd1438 : data_rom <= {16'd4503, 16'd32457};
                15'd1439 : data_rom <= {16'd4506, 16'd32456};
                15'd1440 : data_rom <= {16'd4509, 16'd32456};
                15'd1441 : data_rom <= {16'd4512, 16'd32455};
                15'd1442 : data_rom <= {16'd4515, 16'd32455};
                15'd1443 : data_rom <= {16'd4518, 16'd32454};
                15'd1444 : data_rom <= {16'd4521, 16'd32454};
                15'd1445 : data_rom <= {16'd4525, 16'd32454};
                15'd1446 : data_rom <= {16'd4528, 16'd32453};
                15'd1447 : data_rom <= {16'd4531, 16'd32453};
                15'd1448 : data_rom <= {16'd4534, 16'd32452};
                15'd1449 : data_rom <= {16'd4537, 16'd32452};
                15'd1450 : data_rom <= {16'd4540, 16'd32451};
                15'd1451 : data_rom <= {16'd4543, 16'd32451};
                15'd1452 : data_rom <= {16'd4546, 16'd32451};
                15'd1453 : data_rom <= {16'd4549, 16'd32450};
                15'd1454 : data_rom <= {16'd4553, 16'd32450};
                15'd1455 : data_rom <= {16'd4556, 16'd32449};
                15'd1456 : data_rom <= {16'd4559, 16'd32449};
                15'd1457 : data_rom <= {16'd4562, 16'd32448};
                15'd1458 : data_rom <= {16'd4565, 16'd32448};
                15'd1459 : data_rom <= {16'd4568, 16'd32447};
                15'd1460 : data_rom <= {16'd4571, 16'd32447};
                15'd1461 : data_rom <= {16'd4574, 16'd32447};
                15'd1462 : data_rom <= {16'd4577, 16'd32446};
                15'd1463 : data_rom <= {16'd4581, 16'd32446};
                15'd1464 : data_rom <= {16'd4584, 16'd32445};
                15'd1465 : data_rom <= {16'd4587, 16'd32445};
                15'd1466 : data_rom <= {16'd4590, 16'd32444};
                15'd1467 : data_rom <= {16'd4593, 16'd32444};
                15'd1468 : data_rom <= {16'd4596, 16'd32443};
                15'd1469 : data_rom <= {16'd4599, 16'd32443};
                15'd1470 : data_rom <= {16'd4602, 16'd32443};
                15'd1471 : data_rom <= {16'd4605, 16'd32442};
                15'd1472 : data_rom <= {16'd4609, 16'd32442};
                15'd1473 : data_rom <= {16'd4612, 16'd32441};
                15'd1474 : data_rom <= {16'd4615, 16'd32441};
                15'd1475 : data_rom <= {16'd4618, 16'd32440};
                15'd1476 : data_rom <= {16'd4621, 16'd32440};
                15'd1477 : data_rom <= {16'd4624, 16'd32440};
                15'd1478 : data_rom <= {16'd4627, 16'd32439};
                15'd1479 : data_rom <= {16'd4630, 16'd32439};
                15'd1480 : data_rom <= {16'd4633, 16'd32438};
                15'd1481 : data_rom <= {16'd4637, 16'd32438};
                15'd1482 : data_rom <= {16'd4640, 16'd32437};
                15'd1483 : data_rom <= {16'd4643, 16'd32437};
                15'd1484 : data_rom <= {16'd4646, 16'd32436};
                15'd1485 : data_rom <= {16'd4649, 16'd32436};
                15'd1486 : data_rom <= {16'd4652, 16'd32436};
                15'd1487 : data_rom <= {16'd4655, 16'd32435};
                15'd1488 : data_rom <= {16'd4658, 16'd32435};
                15'd1489 : data_rom <= {16'd4661, 16'd32434};
                15'd1490 : data_rom <= {16'd4665, 16'd32434};
                15'd1491 : data_rom <= {16'd4668, 16'd32433};
                15'd1492 : data_rom <= {16'd4671, 16'd32433};
                15'd1493 : data_rom <= {16'd4674, 16'd32432};
                15'd1494 : data_rom <= {16'd4677, 16'd32432};
                15'd1495 : data_rom <= {16'd4680, 16'd32431};
                15'd1496 : data_rom <= {16'd4683, 16'd32431};
                15'd1497 : data_rom <= {16'd4686, 16'd32431};
                15'd1498 : data_rom <= {16'd4689, 16'd32430};
                15'd1499 : data_rom <= {16'd4693, 16'd32430};
                15'd1500 : data_rom <= {16'd4696, 16'd32429};
                15'd1501 : data_rom <= {16'd4699, 16'd32429};
                15'd1502 : data_rom <= {16'd4702, 16'd32428};
                15'd1503 : data_rom <= {16'd4705, 16'd32428};
                15'd1504 : data_rom <= {16'd4708, 16'd32427};
                15'd1505 : data_rom <= {16'd4711, 16'd32427};
                15'd1506 : data_rom <= {16'd4714, 16'd32427};
                15'd1507 : data_rom <= {16'd4717, 16'd32426};
                15'd1508 : data_rom <= {16'd4721, 16'd32426};
                15'd1509 : data_rom <= {16'd4724, 16'd32425};
                15'd1510 : data_rom <= {16'd4727, 16'd32425};
                15'd1511 : data_rom <= {16'd4730, 16'd32424};
                15'd1512 : data_rom <= {16'd4733, 16'd32424};
                15'd1513 : data_rom <= {16'd4736, 16'd32423};
                15'd1514 : data_rom <= {16'd4739, 16'd32423};
                15'd1515 : data_rom <= {16'd4742, 16'd32422};
                15'd1516 : data_rom <= {16'd4745, 16'd32422};
                15'd1517 : data_rom <= {16'd4749, 16'd32422};
                15'd1518 : data_rom <= {16'd4752, 16'd32421};
                15'd1519 : data_rom <= {16'd4755, 16'd32421};
                15'd1520 : data_rom <= {16'd4758, 16'd32420};
                15'd1521 : data_rom <= {16'd4761, 16'd32420};
                15'd1522 : data_rom <= {16'd4764, 16'd32419};
                15'd1523 : data_rom <= {16'd4767, 16'd32419};
                15'd1524 : data_rom <= {16'd4770, 16'd32418};
                15'd1525 : data_rom <= {16'd4773, 16'd32418};
                15'd1526 : data_rom <= {16'd4776, 16'd32417};
                15'd1527 : data_rom <= {16'd4780, 16'd32417};
                15'd1528 : data_rom <= {16'd4783, 16'd32417};
                15'd1529 : data_rom <= {16'd4786, 16'd32416};
                15'd1530 : data_rom <= {16'd4789, 16'd32416};
                15'd1531 : data_rom <= {16'd4792, 16'd32415};
                15'd1532 : data_rom <= {16'd4795, 16'd32415};
                15'd1533 : data_rom <= {16'd4798, 16'd32414};
                15'd1534 : data_rom <= {16'd4801, 16'd32414};
                15'd1535 : data_rom <= {16'd4804, 16'd32413};
                15'd1536 : data_rom <= {16'd4808, 16'd32413};
                15'd1537 : data_rom <= {16'd4811, 16'd32412};
                15'd1538 : data_rom <= {16'd4814, 16'd32412};
                15'd1539 : data_rom <= {16'd4817, 16'd32411};
                15'd1540 : data_rom <= {16'd4820, 16'd32411};
                15'd1541 : data_rom <= {16'd4823, 16'd32411};
                15'd1542 : data_rom <= {16'd4826, 16'd32410};
                15'd1543 : data_rom <= {16'd4829, 16'd32410};
                15'd1544 : data_rom <= {16'd4832, 16'd32409};
                15'd1545 : data_rom <= {16'd4836, 16'd32409};
                15'd1546 : data_rom <= {16'd4839, 16'd32408};
                15'd1547 : data_rom <= {16'd4842, 16'd32408};
                15'd1548 : data_rom <= {16'd4845, 16'd32407};
                15'd1549 : data_rom <= {16'd4848, 16'd32407};
                15'd1550 : data_rom <= {16'd4851, 16'd32406};
                15'd1551 : data_rom <= {16'd4854, 16'd32406};
                15'd1552 : data_rom <= {16'd4857, 16'd32405};
                15'd1553 : data_rom <= {16'd4860, 16'd32405};
                15'd1554 : data_rom <= {16'd4863, 16'd32404};
                15'd1555 : data_rom <= {16'd4867, 16'd32404};
                15'd1556 : data_rom <= {16'd4870, 16'd32404};
                15'd1557 : data_rom <= {16'd4873, 16'd32403};
                15'd1558 : data_rom <= {16'd4876, 16'd32403};
                15'd1559 : data_rom <= {16'd4879, 16'd32402};
                15'd1560 : data_rom <= {16'd4882, 16'd32402};
                15'd1561 : data_rom <= {16'd4885, 16'd32401};
                15'd1562 : data_rom <= {16'd4888, 16'd32401};
                15'd1563 : data_rom <= {16'd4891, 16'd32400};
                15'd1564 : data_rom <= {16'd4895, 16'd32400};
                15'd1565 : data_rom <= {16'd4898, 16'd32399};
                15'd1566 : data_rom <= {16'd4901, 16'd32399};
                15'd1567 : data_rom <= {16'd4904, 16'd32398};
                15'd1568 : data_rom <= {16'd4907, 16'd32398};
                15'd1569 : data_rom <= {16'd4910, 16'd32397};
                15'd1570 : data_rom <= {16'd4913, 16'd32397};
                15'd1571 : data_rom <= {16'd4916, 16'd32397};
                15'd1572 : data_rom <= {16'd4919, 16'd32396};
                15'd1573 : data_rom <= {16'd4923, 16'd32396};
                15'd1574 : data_rom <= {16'd4926, 16'd32395};
                15'd1575 : data_rom <= {16'd4929, 16'd32395};
                15'd1576 : data_rom <= {16'd4932, 16'd32394};
                15'd1577 : data_rom <= {16'd4935, 16'd32394};
                15'd1578 : data_rom <= {16'd4938, 16'd32393};
                15'd1579 : data_rom <= {16'd4941, 16'd32393};
                15'd1580 : data_rom <= {16'd4944, 16'd32392};
                15'd1581 : data_rom <= {16'd4947, 16'd32392};
                15'd1582 : data_rom <= {16'd4950, 16'd32391};
                15'd1583 : data_rom <= {16'd4954, 16'd32391};
                15'd1584 : data_rom <= {16'd4957, 16'd32390};
                15'd1585 : data_rom <= {16'd4960, 16'd32390};
                15'd1586 : data_rom <= {16'd4963, 16'd32389};
                15'd1587 : data_rom <= {16'd4966, 16'd32389};
                15'd1588 : data_rom <= {16'd4969, 16'd32388};
                15'd1589 : data_rom <= {16'd4972, 16'd32388};
                15'd1590 : data_rom <= {16'd4975, 16'd32388};
                15'd1591 : data_rom <= {16'd4978, 16'd32387};
                15'd1592 : data_rom <= {16'd4982, 16'd32387};
                15'd1593 : data_rom <= {16'd4985, 16'd32386};
                15'd1594 : data_rom <= {16'd4988, 16'd32386};
                15'd1595 : data_rom <= {16'd4991, 16'd32385};
                15'd1596 : data_rom <= {16'd4994, 16'd32385};
                15'd1597 : data_rom <= {16'd4997, 16'd32384};
                15'd1598 : data_rom <= {16'd5000, 16'd32384};
                15'd1599 : data_rom <= {16'd5003, 16'd32383};
                15'd1600 : data_rom <= {16'd5006, 16'd32383};
                15'd1601 : data_rom <= {16'd5009, 16'd32382};
                15'd1602 : data_rom <= {16'd5013, 16'd32382};
                15'd1603 : data_rom <= {16'd5016, 16'd32381};
                15'd1604 : data_rom <= {16'd5019, 16'd32381};
                15'd1605 : data_rom <= {16'd5022, 16'd32380};
                15'd1606 : data_rom <= {16'd5025, 16'd32380};
                15'd1607 : data_rom <= {16'd5028, 16'd32379};
                15'd1608 : data_rom <= {16'd5031, 16'd32379};
                15'd1609 : data_rom <= {16'd5034, 16'd32378};
                15'd1610 : data_rom <= {16'd5037, 16'd32378};
                15'd1611 : data_rom <= {16'd5041, 16'd32377};
                15'd1612 : data_rom <= {16'd5044, 16'd32377};
                15'd1613 : data_rom <= {16'd5047, 16'd32376};
                15'd1614 : data_rom <= {16'd5050, 16'd32376};
                15'd1615 : data_rom <= {16'd5053, 16'd32375};
                15'd1616 : data_rom <= {16'd5056, 16'd32375};
                15'd1617 : data_rom <= {16'd5059, 16'd32375};
                15'd1618 : data_rom <= {16'd5062, 16'd32374};
                15'd1619 : data_rom <= {16'd5065, 16'd32374};
                15'd1620 : data_rom <= {16'd5068, 16'd32373};
                15'd1621 : data_rom <= {16'd5072, 16'd32373};
                15'd1622 : data_rom <= {16'd5075, 16'd32372};
                15'd1623 : data_rom <= {16'd5078, 16'd32372};
                15'd1624 : data_rom <= {16'd5081, 16'd32371};
                15'd1625 : data_rom <= {16'd5084, 16'd32371};
                15'd1626 : data_rom <= {16'd5087, 16'd32370};
                15'd1627 : data_rom <= {16'd5090, 16'd32370};
                15'd1628 : data_rom <= {16'd5093, 16'd32369};
                15'd1629 : data_rom <= {16'd5096, 16'd32369};
                15'd1630 : data_rom <= {16'd5099, 16'd32368};
                15'd1631 : data_rom <= {16'd5103, 16'd32368};
                15'd1632 : data_rom <= {16'd5106, 16'd32367};
                15'd1633 : data_rom <= {16'd5109, 16'd32367};
                15'd1634 : data_rom <= {16'd5112, 16'd32366};
                15'd1635 : data_rom <= {16'd5115, 16'd32366};
                15'd1636 : data_rom <= {16'd5118, 16'd32365};
                15'd1637 : data_rom <= {16'd5121, 16'd32365};
                15'd1638 : data_rom <= {16'd5124, 16'd32364};
                15'd1639 : data_rom <= {16'd5127, 16'd32364};
                15'd1640 : data_rom <= {16'd5131, 16'd32363};
                15'd1641 : data_rom <= {16'd5134, 16'd32363};
                15'd1642 : data_rom <= {16'd5137, 16'd32362};
                15'd1643 : data_rom <= {16'd5140, 16'd32362};
                15'd1644 : data_rom <= {16'd5143, 16'd32361};
                15'd1645 : data_rom <= {16'd5146, 16'd32361};
                15'd1646 : data_rom <= {16'd5149, 16'd32360};
                15'd1647 : data_rom <= {16'd5152, 16'd32360};
                15'd1648 : data_rom <= {16'd5155, 16'd32359};
                15'd1649 : data_rom <= {16'd5158, 16'd32359};
                15'd1650 : data_rom <= {16'd5162, 16'd32358};
                15'd1651 : data_rom <= {16'd5165, 16'd32358};
                15'd1652 : data_rom <= {16'd5168, 16'd32357};
                15'd1653 : data_rom <= {16'd5171, 16'd32357};
                15'd1654 : data_rom <= {16'd5174, 16'd32356};
                15'd1655 : data_rom <= {16'd5177, 16'd32356};
                15'd1656 : data_rom <= {16'd5180, 16'd32355};
                15'd1657 : data_rom <= {16'd5183, 16'd32355};
                15'd1658 : data_rom <= {16'd5186, 16'd32354};
                15'd1659 : data_rom <= {16'd5189, 16'd32354};
                15'd1660 : data_rom <= {16'd5193, 16'd32353};
                15'd1661 : data_rom <= {16'd5196, 16'd32353};
                15'd1662 : data_rom <= {16'd5199, 16'd32352};
                15'd1663 : data_rom <= {16'd5202, 16'd32352};
                15'd1664 : data_rom <= {16'd5205, 16'd32351};
                15'd1665 : data_rom <= {16'd5208, 16'd32351};
                15'd1666 : data_rom <= {16'd5211, 16'd32350};
                15'd1667 : data_rom <= {16'd5214, 16'd32350};
                15'd1668 : data_rom <= {16'd5217, 16'd32349};
                15'd1669 : data_rom <= {16'd5220, 16'd32349};
                15'd1670 : data_rom <= {16'd5224, 16'd32348};
                15'd1671 : data_rom <= {16'd5227, 16'd32348};
                15'd1672 : data_rom <= {16'd5230, 16'd32347};
                15'd1673 : data_rom <= {16'd5233, 16'd32347};
                15'd1674 : data_rom <= {16'd5236, 16'd32346};
                15'd1675 : data_rom <= {16'd5239, 16'd32346};
                15'd1676 : data_rom <= {16'd5242, 16'd32345};
                15'd1677 : data_rom <= {16'd5245, 16'd32345};
                15'd1678 : data_rom <= {16'd5248, 16'd32344};
                15'd1679 : data_rom <= {16'd5251, 16'd32344};
                15'd1680 : data_rom <= {16'd5255, 16'd32343};
                15'd1681 : data_rom <= {16'd5258, 16'd32343};
                15'd1682 : data_rom <= {16'd5261, 16'd32342};
                15'd1683 : data_rom <= {16'd5264, 16'd32342};
                15'd1684 : data_rom <= {16'd5267, 16'd32341};
                15'd1685 : data_rom <= {16'd5270, 16'd32341};
                15'd1686 : data_rom <= {16'd5273, 16'd32340};
                15'd1687 : data_rom <= {16'd5276, 16'd32340};
                15'd1688 : data_rom <= {16'd5279, 16'd32339};
                15'd1689 : data_rom <= {16'd5282, 16'd32339};
                15'd1690 : data_rom <= {16'd5286, 16'd32338};
                15'd1691 : data_rom <= {16'd5289, 16'd32338};
                15'd1692 : data_rom <= {16'd5292, 16'd32337};
                15'd1693 : data_rom <= {16'd5295, 16'd32337};
                15'd1694 : data_rom <= {16'd5298, 16'd32336};
                15'd1695 : data_rom <= {16'd5301, 16'd32336};
                15'd1696 : data_rom <= {16'd5304, 16'd32335};
                15'd1697 : data_rom <= {16'd5307, 16'd32335};
                15'd1698 : data_rom <= {16'd5310, 16'd32334};
                15'd1699 : data_rom <= {16'd5313, 16'd32334};
                15'd1700 : data_rom <= {16'd5317, 16'd32333};
                15'd1701 : data_rom <= {16'd5320, 16'd32333};
                15'd1702 : data_rom <= {16'd5323, 16'd32332};
                15'd1703 : data_rom <= {16'd5326, 16'd32332};
                15'd1704 : data_rom <= {16'd5329, 16'd32331};
                15'd1705 : data_rom <= {16'd5332, 16'd32331};
                15'd1706 : data_rom <= {16'd5335, 16'd32330};
                15'd1707 : data_rom <= {16'd5338, 16'd32330};
                15'd1708 : data_rom <= {16'd5341, 16'd32329};
                15'd1709 : data_rom <= {16'd5344, 16'd32329};
                15'd1710 : data_rom <= {16'd5348, 16'd32328};
                15'd1711 : data_rom <= {16'd5351, 16'd32328};
                15'd1712 : data_rom <= {16'd5354, 16'd32327};
                15'd1713 : data_rom <= {16'd5357, 16'd32327};
                15'd1714 : data_rom <= {16'd5360, 16'd32326};
                15'd1715 : data_rom <= {16'd5363, 16'd32326};
                15'd1716 : data_rom <= {16'd5366, 16'd32325};
                15'd1717 : data_rom <= {16'd5369, 16'd32325};
                15'd1718 : data_rom <= {16'd5372, 16'd32324};
                15'd1719 : data_rom <= {16'd5375, 16'd32323};
                15'd1720 : data_rom <= {16'd5379, 16'd32323};
                15'd1721 : data_rom <= {16'd5382, 16'd32322};
                15'd1722 : data_rom <= {16'd5385, 16'd32322};
                15'd1723 : data_rom <= {16'd5388, 16'd32321};
                15'd1724 : data_rom <= {16'd5391, 16'd32321};
                15'd1725 : data_rom <= {16'd5394, 16'd32320};
                15'd1726 : data_rom <= {16'd5397, 16'd32320};
                15'd1727 : data_rom <= {16'd5400, 16'd32319};
                15'd1728 : data_rom <= {16'd5403, 16'd32319};
                15'd1729 : data_rom <= {16'd5406, 16'd32318};
                15'd1730 : data_rom <= {16'd5410, 16'd32318};
                15'd1731 : data_rom <= {16'd5413, 16'd32317};
                15'd1732 : data_rom <= {16'd5416, 16'd32317};
                15'd1733 : data_rom <= {16'd5419, 16'd32316};
                15'd1734 : data_rom <= {16'd5422, 16'd32316};
                15'd1735 : data_rom <= {16'd5425, 16'd32315};
                15'd1736 : data_rom <= {16'd5428, 16'd32315};
                15'd1737 : data_rom <= {16'd5431, 16'd32314};
                15'd1738 : data_rom <= {16'd5434, 16'd32314};
                15'd1739 : data_rom <= {16'd5437, 16'd32313};
                15'd1740 : data_rom <= {16'd5441, 16'd32313};
                15'd1741 : data_rom <= {16'd5444, 16'd32312};
                15'd1742 : data_rom <= {16'd5447, 16'd32312};
                15'd1743 : data_rom <= {16'd5450, 16'd32311};
                15'd1744 : data_rom <= {16'd5453, 16'd32311};
                15'd1745 : data_rom <= {16'd5456, 16'd32310};
                15'd1746 : data_rom <= {16'd5459, 16'd32309};
                15'd1747 : data_rom <= {16'd5462, 16'd32309};
                15'd1748 : data_rom <= {16'd5465, 16'd32308};
                15'd1749 : data_rom <= {16'd5468, 16'd32308};
                15'd1750 : data_rom <= {16'd5472, 16'd32307};
                15'd1751 : data_rom <= {16'd5475, 16'd32307};
                15'd1752 : data_rom <= {16'd5478, 16'd32306};
                15'd1753 : data_rom <= {16'd5481, 16'd32306};
                15'd1754 : data_rom <= {16'd5484, 16'd32305};
                15'd1755 : data_rom <= {16'd5487, 16'd32305};
                15'd1756 : data_rom <= {16'd5490, 16'd32304};
                15'd1757 : data_rom <= {16'd5493, 16'd32304};
                15'd1758 : data_rom <= {16'd5496, 16'd32303};
                15'd1759 : data_rom <= {16'd5499, 16'd32303};
                15'd1760 : data_rom <= {16'd5502, 16'd32302};
                15'd1761 : data_rom <= {16'd5506, 16'd32302};
                15'd1762 : data_rom <= {16'd5509, 16'd32301};
                15'd1763 : data_rom <= {16'd5512, 16'd32301};
                15'd1764 : data_rom <= {16'd5515, 16'd32300};
                15'd1765 : data_rom <= {16'd5518, 16'd32299};
                15'd1766 : data_rom <= {16'd5521, 16'd32299};
                15'd1767 : data_rom <= {16'd5524, 16'd32298};
                15'd1768 : data_rom <= {16'd5527, 16'd32298};
                15'd1769 : data_rom <= {16'd5530, 16'd32297};
                15'd1770 : data_rom <= {16'd5533, 16'd32297};
                15'd1771 : data_rom <= {16'd5537, 16'd32296};
                15'd1772 : data_rom <= {16'd5540, 16'd32296};
                15'd1773 : data_rom <= {16'd5543, 16'd32295};
                15'd1774 : data_rom <= {16'd5546, 16'd32295};
                15'd1775 : data_rom <= {16'd5549, 16'd32294};
                15'd1776 : data_rom <= {16'd5552, 16'd32294};
                15'd1777 : data_rom <= {16'd5555, 16'd32293};
                15'd1778 : data_rom <= {16'd5558, 16'd32293};
                15'd1779 : data_rom <= {16'd5561, 16'd32292};
                15'd1780 : data_rom <= {16'd5564, 16'd32292};
                15'd1781 : data_rom <= {16'd5568, 16'd32291};
                15'd1782 : data_rom <= {16'd5571, 16'd32290};
                15'd1783 : data_rom <= {16'd5574, 16'd32290};
                15'd1784 : data_rom <= {16'd5577, 16'd32289};
                15'd1785 : data_rom <= {16'd5580, 16'd32289};
                15'd1786 : data_rom <= {16'd5583, 16'd32288};
                15'd1787 : data_rom <= {16'd5586, 16'd32288};
                15'd1788 : data_rom <= {16'd5589, 16'd32287};
                15'd1789 : data_rom <= {16'd5592, 16'd32287};
                15'd1790 : data_rom <= {16'd5595, 16'd32286};
                15'd1791 : data_rom <= {16'd5598, 16'd32286};
                15'd1792 : data_rom <= {16'd5602, 16'd32285};
                15'd1793 : data_rom <= {16'd5605, 16'd32285};
                15'd1794 : data_rom <= {16'd5608, 16'd32284};
                15'd1795 : data_rom <= {16'd5611, 16'd32283};
                15'd1796 : data_rom <= {16'd5614, 16'd32283};
                15'd1797 : data_rom <= {16'd5617, 16'd32282};
                15'd1798 : data_rom <= {16'd5620, 16'd32282};
                15'd1799 : data_rom <= {16'd5623, 16'd32281};
                15'd1800 : data_rom <= {16'd5626, 16'd32281};
                15'd1801 : data_rom <= {16'd5629, 16'd32280};
                15'd1802 : data_rom <= {16'd5633, 16'd32280};
                15'd1803 : data_rom <= {16'd5636, 16'd32279};
                15'd1804 : data_rom <= {16'd5639, 16'd32279};
                15'd1805 : data_rom <= {16'd5642, 16'd32278};
                15'd1806 : data_rom <= {16'd5645, 16'd32278};
                15'd1807 : data_rom <= {16'd5648, 16'd32277};
                15'd1808 : data_rom <= {16'd5651, 16'd32276};
                15'd1809 : data_rom <= {16'd5654, 16'd32276};
                15'd1810 : data_rom <= {16'd5657, 16'd32275};
                15'd1811 : data_rom <= {16'd5660, 16'd32275};
                15'd1812 : data_rom <= {16'd5663, 16'd32274};
                15'd1813 : data_rom <= {16'd5667, 16'd32274};
                15'd1814 : data_rom <= {16'd5670, 16'd32273};
                15'd1815 : data_rom <= {16'd5673, 16'd32273};
                15'd1816 : data_rom <= {16'd5676, 16'd32272};
                15'd1817 : data_rom <= {16'd5679, 16'd32272};
                15'd1818 : data_rom <= {16'd5682, 16'd32271};
                15'd1819 : data_rom <= {16'd5685, 16'd32270};
                15'd1820 : data_rom <= {16'd5688, 16'd32270};
                15'd1821 : data_rom <= {16'd5691, 16'd32269};
                15'd1822 : data_rom <= {16'd5694, 16'd32269};
                15'd1823 : data_rom <= {16'd5698, 16'd32268};
                15'd1824 : data_rom <= {16'd5701, 16'd32268};
                15'd1825 : data_rom <= {16'd5704, 16'd32267};
                15'd1826 : data_rom <= {16'd5707, 16'd32267};
                15'd1827 : data_rom <= {16'd5710, 16'd32266};
                15'd1828 : data_rom <= {16'd5713, 16'd32266};
                15'd1829 : data_rom <= {16'd5716, 16'd32265};
                15'd1830 : data_rom <= {16'd5719, 16'd32264};
                15'd1831 : data_rom <= {16'd5722, 16'd32264};
                15'd1832 : data_rom <= {16'd5725, 16'd32263};
                15'd1833 : data_rom <= {16'd5728, 16'd32263};
                15'd1834 : data_rom <= {16'd5732, 16'd32262};
                15'd1835 : data_rom <= {16'd5735, 16'd32262};
                15'd1836 : data_rom <= {16'd5738, 16'd32261};
                15'd1837 : data_rom <= {16'd5741, 16'd32261};
                15'd1838 : data_rom <= {16'd5744, 16'd32260};
                15'd1839 : data_rom <= {16'd5747, 16'd32260};
                15'd1840 : data_rom <= {16'd5750, 16'd32259};
                15'd1841 : data_rom <= {16'd5753, 16'd32258};
                15'd1842 : data_rom <= {16'd5756, 16'd32258};
                15'd1843 : data_rom <= {16'd5759, 16'd32257};
                15'd1844 : data_rom <= {16'd5762, 16'd32257};
                15'd1845 : data_rom <= {16'd5766, 16'd32256};
                15'd1846 : data_rom <= {16'd5769, 16'd32256};
                15'd1847 : data_rom <= {16'd5772, 16'd32255};
                15'd1848 : data_rom <= {16'd5775, 16'd32255};
                15'd1849 : data_rom <= {16'd5778, 16'd32254};
                15'd1850 : data_rom <= {16'd5781, 16'd32253};
                15'd1851 : data_rom <= {16'd5784, 16'd32253};
                15'd1852 : data_rom <= {16'd5787, 16'd32252};
                15'd1853 : data_rom <= {16'd5790, 16'd32252};
                15'd1854 : data_rom <= {16'd5793, 16'd32251};
                15'd1855 : data_rom <= {16'd5796, 16'd32251};
                15'd1856 : data_rom <= {16'd5800, 16'd32250};
                15'd1857 : data_rom <= {16'd5803, 16'd32250};
                15'd1858 : data_rom <= {16'd5806, 16'd32249};
                15'd1859 : data_rom <= {16'd5809, 16'd32248};
                15'd1860 : data_rom <= {16'd5812, 16'd32248};
                15'd1861 : data_rom <= {16'd5815, 16'd32247};
                15'd1862 : data_rom <= {16'd5818, 16'd32247};
                15'd1863 : data_rom <= {16'd5821, 16'd32246};
                15'd1864 : data_rom <= {16'd5824, 16'd32246};
                15'd1865 : data_rom <= {16'd5827, 16'd32245};
                15'd1866 : data_rom <= {16'd5830, 16'd32245};
                15'd1867 : data_rom <= {16'd5834, 16'd32244};
                15'd1868 : data_rom <= {16'd5837, 16'd32243};
                15'd1869 : data_rom <= {16'd5840, 16'd32243};
                15'd1870 : data_rom <= {16'd5843, 16'd32242};
                15'd1871 : data_rom <= {16'd5846, 16'd32242};
                15'd1872 : data_rom <= {16'd5849, 16'd32241};
                15'd1873 : data_rom <= {16'd5852, 16'd32241};
                15'd1874 : data_rom <= {16'd5855, 16'd32240};
                15'd1875 : data_rom <= {16'd5858, 16'd32239};
                15'd1876 : data_rom <= {16'd5861, 16'd32239};
                15'd1877 : data_rom <= {16'd5864, 16'd32238};
                15'd1878 : data_rom <= {16'd5868, 16'd32238};
                15'd1879 : data_rom <= {16'd5871, 16'd32237};
                15'd1880 : data_rom <= {16'd5874, 16'd32237};
                15'd1881 : data_rom <= {16'd5877, 16'd32236};
                15'd1882 : data_rom <= {16'd5880, 16'd32236};
                15'd1883 : data_rom <= {16'd5883, 16'd32235};
                15'd1884 : data_rom <= {16'd5886, 16'd32234};
                15'd1885 : data_rom <= {16'd5889, 16'd32234};
                15'd1886 : data_rom <= {16'd5892, 16'd32233};
                15'd1887 : data_rom <= {16'd5895, 16'd32233};
                15'd1888 : data_rom <= {16'd5898, 16'd32232};
                15'd1889 : data_rom <= {16'd5902, 16'd32232};
                15'd1890 : data_rom <= {16'd5905, 16'd32231};
                15'd1891 : data_rom <= {16'd5908, 16'd32230};
                15'd1892 : data_rom <= {16'd5911, 16'd32230};
                15'd1893 : data_rom <= {16'd5914, 16'd32229};
                15'd1894 : data_rom <= {16'd5917, 16'd32229};
                15'd1895 : data_rom <= {16'd5920, 16'd32228};
                15'd1896 : data_rom <= {16'd5923, 16'd32228};
                15'd1897 : data_rom <= {16'd5926, 16'd32227};
                15'd1898 : data_rom <= {16'd5929, 16'd32226};
                15'd1899 : data_rom <= {16'd5932, 16'd32226};
                15'd1900 : data_rom <= {16'd5936, 16'd32225};
                15'd1901 : data_rom <= {16'd5939, 16'd32225};
                15'd1902 : data_rom <= {16'd5942, 16'd32224};
                15'd1903 : data_rom <= {16'd5945, 16'd32224};
                15'd1904 : data_rom <= {16'd5948, 16'd32223};
                15'd1905 : data_rom <= {16'd5951, 16'd32222};
                15'd1906 : data_rom <= {16'd5954, 16'd32222};
                15'd1907 : data_rom <= {16'd5957, 16'd32221};
                15'd1908 : data_rom <= {16'd5960, 16'd32221};
                15'd1909 : data_rom <= {16'd5963, 16'd32220};
                15'd1910 : data_rom <= {16'd5966, 16'd32220};
                15'd1911 : data_rom <= {16'd5970, 16'd32219};
                15'd1912 : data_rom <= {16'd5973, 16'd32218};
                15'd1913 : data_rom <= {16'd5976, 16'd32218};
                15'd1914 : data_rom <= {16'd5979, 16'd32217};
                15'd1915 : data_rom <= {16'd5982, 16'd32217};
                15'd1916 : data_rom <= {16'd5985, 16'd32216};
                15'd1917 : data_rom <= {16'd5988, 16'd32216};
                15'd1918 : data_rom <= {16'd5991, 16'd32215};
                15'd1919 : data_rom <= {16'd5994, 16'd32214};
                15'd1920 : data_rom <= {16'd5997, 16'd32214};
                15'd1921 : data_rom <= {16'd6000, 16'd32213};
                15'd1922 : data_rom <= {16'd6004, 16'd32213};
                15'd1923 : data_rom <= {16'd6007, 16'd32212};
                15'd1924 : data_rom <= {16'd6010, 16'd32212};
                15'd1925 : data_rom <= {16'd6013, 16'd32211};
                15'd1926 : data_rom <= {16'd6016, 16'd32210};
                15'd1927 : data_rom <= {16'd6019, 16'd32210};
                15'd1928 : data_rom <= {16'd6022, 16'd32209};
                15'd1929 : data_rom <= {16'd6025, 16'd32209};
                15'd1930 : data_rom <= {16'd6028, 16'd32208};
                15'd1931 : data_rom <= {16'd6031, 16'd32208};
                15'd1932 : data_rom <= {16'd6034, 16'd32207};
                15'd1933 : data_rom <= {16'd6037, 16'd32206};
                15'd1934 : data_rom <= {16'd6041, 16'd32206};
                15'd1935 : data_rom <= {16'd6044, 16'd32205};
                15'd1936 : data_rom <= {16'd6047, 16'd32205};
                15'd1937 : data_rom <= {16'd6050, 16'd32204};
                15'd1938 : data_rom <= {16'd6053, 16'd32204};
                15'd1939 : data_rom <= {16'd6056, 16'd32203};
                15'd1940 : data_rom <= {16'd6059, 16'd32202};
                15'd1941 : data_rom <= {16'd6062, 16'd32202};
                15'd1942 : data_rom <= {16'd6065, 16'd32201};
                15'd1943 : data_rom <= {16'd6068, 16'd32201};
                15'd1944 : data_rom <= {16'd6071, 16'd32200};
                15'd1945 : data_rom <= {16'd6075, 16'd32199};
                15'd1946 : data_rom <= {16'd6078, 16'd32199};
                15'd1947 : data_rom <= {16'd6081, 16'd32198};
                15'd1948 : data_rom <= {16'd6084, 16'd32198};
                15'd1949 : data_rom <= {16'd6087, 16'd32197};
                15'd1950 : data_rom <= {16'd6090, 16'd32197};
                15'd1951 : data_rom <= {16'd6093, 16'd32196};
                15'd1952 : data_rom <= {16'd6096, 16'd32195};
                15'd1953 : data_rom <= {16'd6099, 16'd32195};
                15'd1954 : data_rom <= {16'd6102, 16'd32194};
                15'd1955 : data_rom <= {16'd6105, 16'd32194};
                15'd1956 : data_rom <= {16'd6108, 16'd32193};
                15'd1957 : data_rom <= {16'd6112, 16'd32192};
                15'd1958 : data_rom <= {16'd6115, 16'd32192};
                15'd1959 : data_rom <= {16'd6118, 16'd32191};
                15'd1960 : data_rom <= {16'd6121, 16'd32191};
                15'd1961 : data_rom <= {16'd6124, 16'd32190};
                15'd1962 : data_rom <= {16'd6127, 16'd32189};
                15'd1963 : data_rom <= {16'd6130, 16'd32189};
                15'd1964 : data_rom <= {16'd6133, 16'd32188};
                15'd1965 : data_rom <= {16'd6136, 16'd32188};
                15'd1966 : data_rom <= {16'd6139, 16'd32187};
                15'd1967 : data_rom <= {16'd6142, 16'd32187};
                15'd1968 : data_rom <= {16'd6146, 16'd32186};
                15'd1969 : data_rom <= {16'd6149, 16'd32185};
                15'd1970 : data_rom <= {16'd6152, 16'd32185};
                15'd1971 : data_rom <= {16'd6155, 16'd32184};
                15'd1972 : data_rom <= {16'd6158, 16'd32184};
                15'd1973 : data_rom <= {16'd6161, 16'd32183};
                15'd1974 : data_rom <= {16'd6164, 16'd32182};
                15'd1975 : data_rom <= {16'd6167, 16'd32182};
                15'd1976 : data_rom <= {16'd6170, 16'd32181};
                15'd1977 : data_rom <= {16'd6173, 16'd32181};
                15'd1978 : data_rom <= {16'd6176, 16'd32180};
                15'd1979 : data_rom <= {16'd6179, 16'd32179};
                15'd1980 : data_rom <= {16'd6183, 16'd32179};
                15'd1981 : data_rom <= {16'd6186, 16'd32178};
                15'd1982 : data_rom <= {16'd6189, 16'd32178};
                15'd1983 : data_rom <= {16'd6192, 16'd32177};
                15'd1984 : data_rom <= {16'd6195, 16'd32176};
                15'd1985 : data_rom <= {16'd6198, 16'd32176};
                15'd1986 : data_rom <= {16'd6201, 16'd32175};
                15'd1987 : data_rom <= {16'd6204, 16'd32175};
                15'd1988 : data_rom <= {16'd6207, 16'd32174};
                15'd1989 : data_rom <= {16'd6210, 16'd32174};
                15'd1990 : data_rom <= {16'd6213, 16'd32173};
                15'd1991 : data_rom <= {16'd6216, 16'd32172};
                15'd1992 : data_rom <= {16'd6220, 16'd32172};
                15'd1993 : data_rom <= {16'd6223, 16'd32171};
                15'd1994 : data_rom <= {16'd6226, 16'd32171};
                15'd1995 : data_rom <= {16'd6229, 16'd32170};
                15'd1996 : data_rom <= {16'd6232, 16'd32169};
                15'd1997 : data_rom <= {16'd6235, 16'd32169};
                15'd1998 : data_rom <= {16'd6238, 16'd32168};
                15'd1999 : data_rom <= {16'd6241, 16'd32168};
                15'd2000 : data_rom <= {16'd6244, 16'd32167};
                15'd2001 : data_rom <= {16'd6247, 16'd32166};
                15'd2002 : data_rom <= {16'd6250, 16'd32166};
                15'd2003 : data_rom <= {16'd6253, 16'd32165};
                15'd2004 : data_rom <= {16'd6257, 16'd32165};
                15'd2005 : data_rom <= {16'd6260, 16'd32164};
                15'd2006 : data_rom <= {16'd6263, 16'd32163};
                15'd2007 : data_rom <= {16'd6266, 16'd32163};
                15'd2008 : data_rom <= {16'd6269, 16'd32162};
                15'd2009 : data_rom <= {16'd6272, 16'd32162};
                15'd2010 : data_rom <= {16'd6275, 16'd32161};
                15'd2011 : data_rom <= {16'd6278, 16'd32160};
                15'd2012 : data_rom <= {16'd6281, 16'd32160};
                15'd2013 : data_rom <= {16'd6284, 16'd32159};
                15'd2014 : data_rom <= {16'd6287, 16'd32159};
                15'd2015 : data_rom <= {16'd6291, 16'd32158};
                15'd2016 : data_rom <= {16'd6294, 16'd32157};
                15'd2017 : data_rom <= {16'd6297, 16'd32157};
                15'd2018 : data_rom <= {16'd6300, 16'd32156};
                15'd2019 : data_rom <= {16'd6303, 16'd32156};
                15'd2020 : data_rom <= {16'd6306, 16'd32155};
                15'd2021 : data_rom <= {16'd6309, 16'd32154};
                15'd2022 : data_rom <= {16'd6312, 16'd32154};
                15'd2023 : data_rom <= {16'd6315, 16'd32153};
                15'd2024 : data_rom <= {16'd6318, 16'd32152};
                15'd2025 : data_rom <= {16'd6321, 16'd32152};
                15'd2026 : data_rom <= {16'd6324, 16'd32151};
                15'd2027 : data_rom <= {16'd6327, 16'd32151};
                15'd2028 : data_rom <= {16'd6331, 16'd32150};
                15'd2029 : data_rom <= {16'd6334, 16'd32149};
                15'd2030 : data_rom <= {16'd6337, 16'd32149};
                15'd2031 : data_rom <= {16'd6340, 16'd32148};
                15'd2032 : data_rom <= {16'd6343, 16'd32148};
                15'd2033 : data_rom <= {16'd6346, 16'd32147};
                15'd2034 : data_rom <= {16'd6349, 16'd32146};
                15'd2035 : data_rom <= {16'd6352, 16'd32146};
                15'd2036 : data_rom <= {16'd6355, 16'd32145};
                15'd2037 : data_rom <= {16'd6358, 16'd32145};
                15'd2038 : data_rom <= {16'd6361, 16'd32144};
                15'd2039 : data_rom <= {16'd6364, 16'd32143};
                15'd2040 : data_rom <= {16'd6368, 16'd32143};
                15'd2041 : data_rom <= {16'd6371, 16'd32142};
                15'd2042 : data_rom <= {16'd6374, 16'd32142};
                15'd2043 : data_rom <= {16'd6377, 16'd32141};
                15'd2044 : data_rom <= {16'd6380, 16'd32140};
                15'd2045 : data_rom <= {16'd6383, 16'd32140};
                15'd2046 : data_rom <= {16'd6386, 16'd32139};
                15'd2047 : data_rom <= {16'd6389, 16'd32138};
                15'd2048 : data_rom <= {16'd6392, 16'd32138};
                15'd2049 : data_rom <= {16'd6395, 16'd32137};
                15'd2050 : data_rom <= {16'd6398, 16'd32137};
                15'd2051 : data_rom <= {16'd6401, 16'd32136};
                15'd2052 : data_rom <= {16'd6405, 16'd32135};
                15'd2053 : data_rom <= {16'd6408, 16'd32135};
                15'd2054 : data_rom <= {16'd6411, 16'd32134};
                15'd2055 : data_rom <= {16'd6414, 16'd32134};
                15'd2056 : data_rom <= {16'd6417, 16'd32133};
                15'd2057 : data_rom <= {16'd6420, 16'd32132};
                15'd2058 : data_rom <= {16'd6423, 16'd32132};
                15'd2059 : data_rom <= {16'd6426, 16'd32131};
                15'd2060 : data_rom <= {16'd6429, 16'd32130};
                15'd2061 : data_rom <= {16'd6432, 16'd32130};
                15'd2062 : data_rom <= {16'd6435, 16'd32129};
                15'd2063 : data_rom <= {16'd6438, 16'd32129};
                15'd2064 : data_rom <= {16'd6442, 16'd32128};
                15'd2065 : data_rom <= {16'd6445, 16'd32127};
                15'd2066 : data_rom <= {16'd6448, 16'd32127};
                15'd2067 : data_rom <= {16'd6451, 16'd32126};
                15'd2068 : data_rom <= {16'd6454, 16'd32126};
                15'd2069 : data_rom <= {16'd6457, 16'd32125};
                15'd2070 : data_rom <= {16'd6460, 16'd32124};
                15'd2071 : data_rom <= {16'd6463, 16'd32124};
                15'd2072 : data_rom <= {16'd6466, 16'd32123};
                15'd2073 : data_rom <= {16'd6469, 16'd32122};
                15'd2074 : data_rom <= {16'd6472, 16'd32122};
                15'd2075 : data_rom <= {16'd6475, 16'd32121};
                15'd2076 : data_rom <= {16'd6478, 16'd32121};
                15'd2077 : data_rom <= {16'd6482, 16'd32120};
                15'd2078 : data_rom <= {16'd6485, 16'd32119};
                15'd2079 : data_rom <= {16'd6488, 16'd32119};
                15'd2080 : data_rom <= {16'd6491, 16'd32118};
                15'd2081 : data_rom <= {16'd6494, 16'd32117};
                15'd2082 : data_rom <= {16'd6497, 16'd32117};
                15'd2083 : data_rom <= {16'd6500, 16'd32116};
                15'd2084 : data_rom <= {16'd6503, 16'd32116};
                15'd2085 : data_rom <= {16'd6506, 16'd32115};
                15'd2086 : data_rom <= {16'd6509, 16'd32114};
                15'd2087 : data_rom <= {16'd6512, 16'd32114};
                15'd2088 : data_rom <= {16'd6515, 16'd32113};
                15'd2089 : data_rom <= {16'd6518, 16'd32112};
                15'd2090 : data_rom <= {16'd6522, 16'd32112};
                15'd2091 : data_rom <= {16'd6525, 16'd32111};
                15'd2092 : data_rom <= {16'd6528, 16'd32111};
                15'd2093 : data_rom <= {16'd6531, 16'd32110};
                15'd2094 : data_rom <= {16'd6534, 16'd32109};
                15'd2095 : data_rom <= {16'd6537, 16'd32109};
                15'd2096 : data_rom <= {16'd6540, 16'd32108};
                15'd2097 : data_rom <= {16'd6543, 16'd32107};
                15'd2098 : data_rom <= {16'd6546, 16'd32107};
                15'd2099 : data_rom <= {16'd6549, 16'd32106};
                15'd2100 : data_rom <= {16'd6552, 16'd32106};
                15'd2101 : data_rom <= {16'd6555, 16'd32105};
                15'd2102 : data_rom <= {16'd6559, 16'd32104};
                15'd2103 : data_rom <= {16'd6562, 16'd32104};
                15'd2104 : data_rom <= {16'd6565, 16'd32103};
                15'd2105 : data_rom <= {16'd6568, 16'd32102};
                15'd2106 : data_rom <= {16'd6571, 16'd32102};
                15'd2107 : data_rom <= {16'd6574, 16'd32101};
                15'd2108 : data_rom <= {16'd6577, 16'd32101};
                15'd2109 : data_rom <= {16'd6580, 16'd32100};
                15'd2110 : data_rom <= {16'd6583, 16'd32099};
                15'd2111 : data_rom <= {16'd6586, 16'd32099};
                15'd2112 : data_rom <= {16'd6589, 16'd32098};
                15'd2113 : data_rom <= {16'd6592, 16'd32097};
                15'd2114 : data_rom <= {16'd6595, 16'd32097};
                15'd2115 : data_rom <= {16'd6599, 16'd32096};
                15'd2116 : data_rom <= {16'd6602, 16'd32096};
                15'd2117 : data_rom <= {16'd6605, 16'd32095};
                15'd2118 : data_rom <= {16'd6608, 16'd32094};
                15'd2119 : data_rom <= {16'd6611, 16'd32094};
                15'd2120 : data_rom <= {16'd6614, 16'd32093};
                15'd2121 : data_rom <= {16'd6617, 16'd32092};
                15'd2122 : data_rom <= {16'd6620, 16'd32092};
                15'd2123 : data_rom <= {16'd6623, 16'd32091};
                15'd2124 : data_rom <= {16'd6626, 16'd32090};
                15'd2125 : data_rom <= {16'd6629, 16'd32090};
                15'd2126 : data_rom <= {16'd6632, 16'd32089};
                15'd2127 : data_rom <= {16'd6635, 16'd32089};
                15'd2128 : data_rom <= {16'd6639, 16'd32088};
                15'd2129 : data_rom <= {16'd6642, 16'd32087};
                15'd2130 : data_rom <= {16'd6645, 16'd32087};
                15'd2131 : data_rom <= {16'd6648, 16'd32086};
                15'd2132 : data_rom <= {16'd6651, 16'd32085};
                15'd2133 : data_rom <= {16'd6654, 16'd32085};
                15'd2134 : data_rom <= {16'd6657, 16'd32084};
                15'd2135 : data_rom <= {16'd6660, 16'd32083};
                15'd2136 : data_rom <= {16'd6663, 16'd32083};
                15'd2137 : data_rom <= {16'd6666, 16'd32082};
                15'd2138 : data_rom <= {16'd6669, 16'd32082};
                15'd2139 : data_rom <= {16'd6672, 16'd32081};
                15'd2140 : data_rom <= {16'd6675, 16'd32080};
                15'd2141 : data_rom <= {16'd6679, 16'd32080};
                15'd2142 : data_rom <= {16'd6682, 16'd32079};
                15'd2143 : data_rom <= {16'd6685, 16'd32078};
                15'd2144 : data_rom <= {16'd6688, 16'd32078};
                15'd2145 : data_rom <= {16'd6691, 16'd32077};
                15'd2146 : data_rom <= {16'd6694, 16'd32076};
                15'd2147 : data_rom <= {16'd6697, 16'd32076};
                15'd2148 : data_rom <= {16'd6700, 16'd32075};
                15'd2149 : data_rom <= {16'd6703, 16'd32074};
                15'd2150 : data_rom <= {16'd6706, 16'd32074};
                15'd2151 : data_rom <= {16'd6709, 16'd32073};
                15'd2152 : data_rom <= {16'd6712, 16'd32073};
                15'd2153 : data_rom <= {16'd6715, 16'd32072};
                15'd2154 : data_rom <= {16'd6718, 16'd32071};
                15'd2155 : data_rom <= {16'd6722, 16'd32071};
                15'd2156 : data_rom <= {16'd6725, 16'd32070};
                15'd2157 : data_rom <= {16'd6728, 16'd32069};
                15'd2158 : data_rom <= {16'd6731, 16'd32069};
                15'd2159 : data_rom <= {16'd6734, 16'd32068};
                15'd2160 : data_rom <= {16'd6737, 16'd32067};
                15'd2161 : data_rom <= {16'd6740, 16'd32067};
                15'd2162 : data_rom <= {16'd6743, 16'd32066};
                15'd2163 : data_rom <= {16'd6746, 16'd32065};
                15'd2164 : data_rom <= {16'd6749, 16'd32065};
                15'd2165 : data_rom <= {16'd6752, 16'd32064};
                15'd2166 : data_rom <= {16'd6755, 16'd32063};
                15'd2167 : data_rom <= {16'd6758, 16'd32063};
                15'd2168 : data_rom <= {16'd6762, 16'd32062};
                15'd2169 : data_rom <= {16'd6765, 16'd32062};
                15'd2170 : data_rom <= {16'd6768, 16'd32061};
                15'd2171 : data_rom <= {16'd6771, 16'd32060};
                15'd2172 : data_rom <= {16'd6774, 16'd32060};
                15'd2173 : data_rom <= {16'd6777, 16'd32059};
                15'd2174 : data_rom <= {16'd6780, 16'd32058};
                15'd2175 : data_rom <= {16'd6783, 16'd32058};
                15'd2176 : data_rom <= {16'd6786, 16'd32057};
                15'd2177 : data_rom <= {16'd6789, 16'd32056};
                15'd2178 : data_rom <= {16'd6792, 16'd32056};
                15'd2179 : data_rom <= {16'd6795, 16'd32055};
                15'd2180 : data_rom <= {16'd6798, 16'd32054};
                15'd2181 : data_rom <= {16'd6801, 16'd32054};
                15'd2182 : data_rom <= {16'd6805, 16'd32053};
                15'd2183 : data_rom <= {16'd6808, 16'd32052};
                15'd2184 : data_rom <= {16'd6811, 16'd32052};
                15'd2185 : data_rom <= {16'd6814, 16'd32051};
                15'd2186 : data_rom <= {16'd6817, 16'd32050};
                15'd2187 : data_rom <= {16'd6820, 16'd32050};
                15'd2188 : data_rom <= {16'd6823, 16'd32049};
                15'd2189 : data_rom <= {16'd6826, 16'd32049};
                15'd2190 : data_rom <= {16'd6829, 16'd32048};
                15'd2191 : data_rom <= {16'd6832, 16'd32047};
                15'd2192 : data_rom <= {16'd6835, 16'd32047};
                15'd2193 : data_rom <= {16'd6838, 16'd32046};
                15'd2194 : data_rom <= {16'd6841, 16'd32045};
                15'd2195 : data_rom <= {16'd6845, 16'd32045};
                15'd2196 : data_rom <= {16'd6848, 16'd32044};
                15'd2197 : data_rom <= {16'd6851, 16'd32043};
                15'd2198 : data_rom <= {16'd6854, 16'd32043};
                15'd2199 : data_rom <= {16'd6857, 16'd32042};
                15'd2200 : data_rom <= {16'd6860, 16'd32041};
                15'd2201 : data_rom <= {16'd6863, 16'd32041};
                15'd2202 : data_rom <= {16'd6866, 16'd32040};
                15'd2203 : data_rom <= {16'd6869, 16'd32039};
                15'd2204 : data_rom <= {16'd6872, 16'd32039};
                15'd2205 : data_rom <= {16'd6875, 16'd32038};
                15'd2206 : data_rom <= {16'd6878, 16'd32037};
                15'd2207 : data_rom <= {16'd6881, 16'd32037};
                15'd2208 : data_rom <= {16'd6884, 16'd32036};
                15'd2209 : data_rom <= {16'd6888, 16'd32035};
                15'd2210 : data_rom <= {16'd6891, 16'd32035};
                15'd2211 : data_rom <= {16'd6894, 16'd32034};
                15'd2212 : data_rom <= {16'd6897, 16'd32033};
                15'd2213 : data_rom <= {16'd6900, 16'd32033};
                15'd2214 : data_rom <= {16'd6903, 16'd32032};
                15'd2215 : data_rom <= {16'd6906, 16'd32031};
                15'd2216 : data_rom <= {16'd6909, 16'd32031};
                15'd2217 : data_rom <= {16'd6912, 16'd32030};
                15'd2218 : data_rom <= {16'd6915, 16'd32029};
                15'd2219 : data_rom <= {16'd6918, 16'd32029};
                15'd2220 : data_rom <= {16'd6921, 16'd32028};
                15'd2221 : data_rom <= {16'd6924, 16'd32027};
                15'd2222 : data_rom <= {16'd6927, 16'd32027};
                15'd2223 : data_rom <= {16'd6931, 16'd32026};
                15'd2224 : data_rom <= {16'd6934, 16'd32025};
                15'd2225 : data_rom <= {16'd6937, 16'd32025};
                15'd2226 : data_rom <= {16'd6940, 16'd32024};
                15'd2227 : data_rom <= {16'd6943, 16'd32023};
                15'd2228 : data_rom <= {16'd6946, 16'd32023};
                15'd2229 : data_rom <= {16'd6949, 16'd32022};
                15'd2230 : data_rom <= {16'd6952, 16'd32021};
                15'd2231 : data_rom <= {16'd6955, 16'd32021};
                15'd2232 : data_rom <= {16'd6958, 16'd32020};
                15'd2233 : data_rom <= {16'd6961, 16'd32019};
                15'd2234 : data_rom <= {16'd6964, 16'd32019};
                15'd2235 : data_rom <= {16'd6967, 16'd32018};
                15'd2236 : data_rom <= {16'd6970, 16'd32017};
                15'd2237 : data_rom <= {16'd6973, 16'd32017};
                15'd2238 : data_rom <= {16'd6977, 16'd32016};
                15'd2239 : data_rom <= {16'd6980, 16'd32015};
                15'd2240 : data_rom <= {16'd6983, 16'd32015};
                15'd2241 : data_rom <= {16'd6986, 16'd32014};
                15'd2242 : data_rom <= {16'd6989, 16'd32013};
                15'd2243 : data_rom <= {16'd6992, 16'd32013};
                15'd2244 : data_rom <= {16'd6995, 16'd32012};
                15'd2245 : data_rom <= {16'd6998, 16'd32011};
                15'd2246 : data_rom <= {16'd7001, 16'd32011};
                15'd2247 : data_rom <= {16'd7004, 16'd32010};
                15'd2248 : data_rom <= {16'd7007, 16'd32009};
                15'd2249 : data_rom <= {16'd7010, 16'd32009};
                15'd2250 : data_rom <= {16'd7013, 16'd32008};
                15'd2251 : data_rom <= {16'd7016, 16'd32007};
                15'd2252 : data_rom <= {16'd7020, 16'd32007};
                15'd2253 : data_rom <= {16'd7023, 16'd32006};
                15'd2254 : data_rom <= {16'd7026, 16'd32005};
                15'd2255 : data_rom <= {16'd7029, 16'd32005};
                15'd2256 : data_rom <= {16'd7032, 16'd32004};
                15'd2257 : data_rom <= {16'd7035, 16'd32003};
                15'd2258 : data_rom <= {16'd7038, 16'd32003};
                15'd2259 : data_rom <= {16'd7041, 16'd32002};
                15'd2260 : data_rom <= {16'd7044, 16'd32001};
                15'd2261 : data_rom <= {16'd7047, 16'd32001};
                15'd2262 : data_rom <= {16'd7050, 16'd32000};
                15'd2263 : data_rom <= {16'd7053, 16'd31999};
                15'd2264 : data_rom <= {16'd7056, 16'd31999};
                15'd2265 : data_rom <= {16'd7059, 16'd31998};
                15'd2266 : data_rom <= {16'd7062, 16'd31997};
                15'd2267 : data_rom <= {16'd7066, 16'd31997};
                15'd2268 : data_rom <= {16'd7069, 16'd31996};
                15'd2269 : data_rom <= {16'd7072, 16'd31995};
                15'd2270 : data_rom <= {16'd7075, 16'd31995};
                15'd2271 : data_rom <= {16'd7078, 16'd31994};
                15'd2272 : data_rom <= {16'd7081, 16'd31993};
                15'd2273 : data_rom <= {16'd7084, 16'd31993};
                15'd2274 : data_rom <= {16'd7087, 16'd31992};
                15'd2275 : data_rom <= {16'd7090, 16'd31991};
                15'd2276 : data_rom <= {16'd7093, 16'd31990};
                15'd2277 : data_rom <= {16'd7096, 16'd31990};
                15'd2278 : data_rom <= {16'd7099, 16'd31989};
                15'd2279 : data_rom <= {16'd7102, 16'd31988};
                15'd2280 : data_rom <= {16'd7105, 16'd31988};
                15'd2281 : data_rom <= {16'd7108, 16'd31987};
                15'd2282 : data_rom <= {16'd7112, 16'd31986};
                15'd2283 : data_rom <= {16'd7115, 16'd31986};
                15'd2284 : data_rom <= {16'd7118, 16'd31985};
                15'd2285 : data_rom <= {16'd7121, 16'd31984};
                15'd2286 : data_rom <= {16'd7124, 16'd31984};
                15'd2287 : data_rom <= {16'd7127, 16'd31983};
                15'd2288 : data_rom <= {16'd7130, 16'd31982};
                15'd2289 : data_rom <= {16'd7133, 16'd31982};
                15'd2290 : data_rom <= {16'd7136, 16'd31981};
                15'd2291 : data_rom <= {16'd7139, 16'd31980};
                15'd2292 : data_rom <= {16'd7142, 16'd31980};
                15'd2293 : data_rom <= {16'd7145, 16'd31979};
                15'd2294 : data_rom <= {16'd7148, 16'd31978};
                15'd2295 : data_rom <= {16'd7151, 16'd31977};
                15'd2296 : data_rom <= {16'd7154, 16'd31977};
                15'd2297 : data_rom <= {16'd7158, 16'd31976};
                15'd2298 : data_rom <= {16'd7161, 16'd31975};
                15'd2299 : data_rom <= {16'd7164, 16'd31975};
                15'd2300 : data_rom <= {16'd7167, 16'd31974};
                15'd2301 : data_rom <= {16'd7170, 16'd31973};
                15'd2302 : data_rom <= {16'd7173, 16'd31973};
                15'd2303 : data_rom <= {16'd7176, 16'd31972};
                15'd2304 : data_rom <= {16'd7179, 16'd31971};
                15'd2305 : data_rom <= {16'd7182, 16'd31971};
                15'd2306 : data_rom <= {16'd7185, 16'd31970};
                15'd2307 : data_rom <= {16'd7188, 16'd31969};
                15'd2308 : data_rom <= {16'd7191, 16'd31969};
                15'd2309 : data_rom <= {16'd7194, 16'd31968};
                15'd2310 : data_rom <= {16'd7197, 16'd31967};
                15'd2311 : data_rom <= {16'd7200, 16'd31966};
                15'd2312 : data_rom <= {16'd7204, 16'd31966};
                15'd2313 : data_rom <= {16'd7207, 16'd31965};
                15'd2314 : data_rom <= {16'd7210, 16'd31964};
                15'd2315 : data_rom <= {16'd7213, 16'd31964};
                15'd2316 : data_rom <= {16'd7216, 16'd31963};
                15'd2317 : data_rom <= {16'd7219, 16'd31962};
                15'd2318 : data_rom <= {16'd7222, 16'd31962};
                15'd2319 : data_rom <= {16'd7225, 16'd31961};
                15'd2320 : data_rom <= {16'd7228, 16'd31960};
                15'd2321 : data_rom <= {16'd7231, 16'd31960};
                15'd2322 : data_rom <= {16'd7234, 16'd31959};
                15'd2323 : data_rom <= {16'd7237, 16'd31958};
                15'd2324 : data_rom <= {16'd7240, 16'd31957};
                15'd2325 : data_rom <= {16'd7243, 16'd31957};
                15'd2326 : data_rom <= {16'd7246, 16'd31956};
                15'd2327 : data_rom <= {16'd7249, 16'd31955};
                15'd2328 : data_rom <= {16'd7253, 16'd31955};
                15'd2329 : data_rom <= {16'd7256, 16'd31954};
                15'd2330 : data_rom <= {16'd7259, 16'd31953};
                15'd2331 : data_rom <= {16'd7262, 16'd31953};
                15'd2332 : data_rom <= {16'd7265, 16'd31952};
                15'd2333 : data_rom <= {16'd7268, 16'd31951};
                15'd2334 : data_rom <= {16'd7271, 16'd31951};
                15'd2335 : data_rom <= {16'd7274, 16'd31950};
                15'd2336 : data_rom <= {16'd7277, 16'd31949};
                15'd2337 : data_rom <= {16'd7280, 16'd31948};
                15'd2338 : data_rom <= {16'd7283, 16'd31948};
                15'd2339 : data_rom <= {16'd7286, 16'd31947};
                15'd2340 : data_rom <= {16'd7289, 16'd31946};
                15'd2341 : data_rom <= {16'd7292, 16'd31946};
                15'd2342 : data_rom <= {16'd7295, 16'd31945};
                15'd2343 : data_rom <= {16'd7298, 16'd31944};
                15'd2344 : data_rom <= {16'd7302, 16'd31944};
                15'd2345 : data_rom <= {16'd7305, 16'd31943};
                15'd2346 : data_rom <= {16'd7308, 16'd31942};
                15'd2347 : data_rom <= {16'd7311, 16'd31941};
                15'd2348 : data_rom <= {16'd7314, 16'd31941};
                15'd2349 : data_rom <= {16'd7317, 16'd31940};
                15'd2350 : data_rom <= {16'd7320, 16'd31939};
                15'd2351 : data_rom <= {16'd7323, 16'd31939};
                15'd2352 : data_rom <= {16'd7326, 16'd31938};
                15'd2353 : data_rom <= {16'd7329, 16'd31937};
                15'd2354 : data_rom <= {16'd7332, 16'd31937};
                15'd2355 : data_rom <= {16'd7335, 16'd31936};
                15'd2356 : data_rom <= {16'd7338, 16'd31935};
                15'd2357 : data_rom <= {16'd7341, 16'd31934};
                15'd2358 : data_rom <= {16'd7344, 16'd31934};
                15'd2359 : data_rom <= {16'd7347, 16'd31933};
                15'd2360 : data_rom <= {16'd7351, 16'd31932};
                15'd2361 : data_rom <= {16'd7354, 16'd31932};
                15'd2362 : data_rom <= {16'd7357, 16'd31931};
                15'd2363 : data_rom <= {16'd7360, 16'd31930};
                15'd2364 : data_rom <= {16'd7363, 16'd31929};
                15'd2365 : data_rom <= {16'd7366, 16'd31929};
                15'd2366 : data_rom <= {16'd7369, 16'd31928};
                15'd2367 : data_rom <= {16'd7372, 16'd31927};
                15'd2368 : data_rom <= {16'd7375, 16'd31927};
                15'd2369 : data_rom <= {16'd7378, 16'd31926};
                15'd2370 : data_rom <= {16'd7381, 16'd31925};
                15'd2371 : data_rom <= {16'd7384, 16'd31925};
                15'd2372 : data_rom <= {16'd7387, 16'd31924};
                15'd2373 : data_rom <= {16'd7390, 16'd31923};
                15'd2374 : data_rom <= {16'd7393, 16'd31922};
                15'd2375 : data_rom <= {16'd7396, 16'd31922};
                15'd2376 : data_rom <= {16'd7400, 16'd31921};
                15'd2377 : data_rom <= {16'd7403, 16'd31920};
                15'd2378 : data_rom <= {16'd7406, 16'd31920};
                15'd2379 : data_rom <= {16'd7409, 16'd31919};
                15'd2380 : data_rom <= {16'd7412, 16'd31918};
                15'd2381 : data_rom <= {16'd7415, 16'd31917};
                15'd2382 : data_rom <= {16'd7418, 16'd31917};
                15'd2383 : data_rom <= {16'd7421, 16'd31916};
                15'd2384 : data_rom <= {16'd7424, 16'd31915};
                15'd2385 : data_rom <= {16'd7427, 16'd31915};
                15'd2386 : data_rom <= {16'd7430, 16'd31914};
                15'd2387 : data_rom <= {16'd7433, 16'd31913};
                15'd2388 : data_rom <= {16'd7436, 16'd31912};
                15'd2389 : data_rom <= {16'd7439, 16'd31912};
                15'd2390 : data_rom <= {16'd7442, 16'd31911};
                15'd2391 : data_rom <= {16'd7445, 16'd31910};
                15'd2392 : data_rom <= {16'd7448, 16'd31910};
                15'd2393 : data_rom <= {16'd7452, 16'd31909};
                15'd2394 : data_rom <= {16'd7455, 16'd31908};
                15'd2395 : data_rom <= {16'd7458, 16'd31907};
                15'd2396 : data_rom <= {16'd7461, 16'd31907};
                15'd2397 : data_rom <= {16'd7464, 16'd31906};
                15'd2398 : data_rom <= {16'd7467, 16'd31905};
                15'd2399 : data_rom <= {16'd7470, 16'd31905};
                15'd2400 : data_rom <= {16'd7473, 16'd31904};
                15'd2401 : data_rom <= {16'd7476, 16'd31903};
                15'd2402 : data_rom <= {16'd7479, 16'd31902};
                15'd2403 : data_rom <= {16'd7482, 16'd31902};
                15'd2404 : data_rom <= {16'd7485, 16'd31901};
                15'd2405 : data_rom <= {16'd7488, 16'd31900};
                15'd2406 : data_rom <= {16'd7491, 16'd31900};
                15'd2407 : data_rom <= {16'd7494, 16'd31899};
                15'd2408 : data_rom <= {16'd7497, 16'd31898};
                15'd2409 : data_rom <= {16'd7500, 16'd31897};
                15'd2410 : data_rom <= {16'd7504, 16'd31897};
                15'd2411 : data_rom <= {16'd7507, 16'd31896};
                15'd2412 : data_rom <= {16'd7510, 16'd31895};
                15'd2413 : data_rom <= {16'd7513, 16'd31895};
                15'd2414 : data_rom <= {16'd7516, 16'd31894};
                15'd2415 : data_rom <= {16'd7519, 16'd31893};
                15'd2416 : data_rom <= {16'd7522, 16'd31892};
                15'd2417 : data_rom <= {16'd7525, 16'd31892};
                15'd2418 : data_rom <= {16'd7528, 16'd31891};
                15'd2419 : data_rom <= {16'd7531, 16'd31890};
                15'd2420 : data_rom <= {16'd7534, 16'd31889};
                15'd2421 : data_rom <= {16'd7537, 16'd31889};
                15'd2422 : data_rom <= {16'd7540, 16'd31888};
                15'd2423 : data_rom <= {16'd7543, 16'd31887};
                15'd2424 : data_rom <= {16'd7546, 16'd31887};
                15'd2425 : data_rom <= {16'd7549, 16'd31886};
                15'd2426 : data_rom <= {16'd7552, 16'd31885};
                15'd2427 : data_rom <= {16'd7556, 16'd31884};
                15'd2428 : data_rom <= {16'd7559, 16'd31884};
                15'd2429 : data_rom <= {16'd7562, 16'd31883};
                15'd2430 : data_rom <= {16'd7565, 16'd31882};
                15'd2431 : data_rom <= {16'd7568, 16'd31882};
                15'd2432 : data_rom <= {16'd7571, 16'd31881};
                15'd2433 : data_rom <= {16'd7574, 16'd31880};
                15'd2434 : data_rom <= {16'd7577, 16'd31879};
                15'd2435 : data_rom <= {16'd7580, 16'd31879};
                15'd2436 : data_rom <= {16'd7583, 16'd31878};
                15'd2437 : data_rom <= {16'd7586, 16'd31877};
                15'd2438 : data_rom <= {16'd7589, 16'd31876};
                15'd2439 : data_rom <= {16'd7592, 16'd31876};
                15'd2440 : data_rom <= {16'd7595, 16'd31875};
                15'd2441 : data_rom <= {16'd7598, 16'd31874};
                15'd2442 : data_rom <= {16'd7601, 16'd31874};
                15'd2443 : data_rom <= {16'd7604, 16'd31873};
                15'd2444 : data_rom <= {16'd7607, 16'd31872};
                15'd2445 : data_rom <= {16'd7611, 16'd31871};
                15'd2446 : data_rom <= {16'd7614, 16'd31871};
                15'd2447 : data_rom <= {16'd7617, 16'd31870};
                15'd2448 : data_rom <= {16'd7620, 16'd31869};
                15'd2449 : data_rom <= {16'd7623, 16'd31868};
                15'd2450 : data_rom <= {16'd7626, 16'd31868};
                15'd2451 : data_rom <= {16'd7629, 16'd31867};
                15'd2452 : data_rom <= {16'd7632, 16'd31866};
                15'd2453 : data_rom <= {16'd7635, 16'd31865};
                15'd2454 : data_rom <= {16'd7638, 16'd31865};
                15'd2455 : data_rom <= {16'd7641, 16'd31864};
                15'd2456 : data_rom <= {16'd7644, 16'd31863};
                15'd2457 : data_rom <= {16'd7647, 16'd31863};
                15'd2458 : data_rom <= {16'd7650, 16'd31862};
                15'd2459 : data_rom <= {16'd7653, 16'd31861};
                15'd2460 : data_rom <= {16'd7656, 16'd31860};
                15'd2461 : data_rom <= {16'd7659, 16'd31860};
                15'd2462 : data_rom <= {16'd7662, 16'd31859};
                15'd2463 : data_rom <= {16'd7666, 16'd31858};
                15'd2464 : data_rom <= {16'd7669, 16'd31857};
                15'd2465 : data_rom <= {16'd7672, 16'd31857};
                15'd2466 : data_rom <= {16'd7675, 16'd31856};
                15'd2467 : data_rom <= {16'd7678, 16'd31855};
                15'd2468 : data_rom <= {16'd7681, 16'd31854};
                15'd2469 : data_rom <= {16'd7684, 16'd31854};
                15'd2470 : data_rom <= {16'd7687, 16'd31853};
                15'd2471 : data_rom <= {16'd7690, 16'd31852};
                15'd2472 : data_rom <= {16'd7693, 16'd31852};
                15'd2473 : data_rom <= {16'd7696, 16'd31851};
                15'd2474 : data_rom <= {16'd7699, 16'd31850};
                15'd2475 : data_rom <= {16'd7702, 16'd31849};
                15'd2476 : data_rom <= {16'd7705, 16'd31849};
                15'd2477 : data_rom <= {16'd7708, 16'd31848};
                15'd2478 : data_rom <= {16'd7711, 16'd31847};
                15'd2479 : data_rom <= {16'd7714, 16'd31846};
                15'd2480 : data_rom <= {16'd7717, 16'd31846};
                15'd2481 : data_rom <= {16'd7720, 16'd31845};
                15'd2482 : data_rom <= {16'd7724, 16'd31844};
                15'd2483 : data_rom <= {16'd7727, 16'd31843};
                15'd2484 : data_rom <= {16'd7730, 16'd31843};
                15'd2485 : data_rom <= {16'd7733, 16'd31842};
                15'd2486 : data_rom <= {16'd7736, 16'd31841};
                15'd2487 : data_rom <= {16'd7739, 16'd31840};
                15'd2488 : data_rom <= {16'd7742, 16'd31840};
                15'd2489 : data_rom <= {16'd7745, 16'd31839};
                15'd2490 : data_rom <= {16'd7748, 16'd31838};
                15'd2491 : data_rom <= {16'd7751, 16'd31837};
                15'd2492 : data_rom <= {16'd7754, 16'd31837};
                15'd2493 : data_rom <= {16'd7757, 16'd31836};
                15'd2494 : data_rom <= {16'd7760, 16'd31835};
                15'd2495 : data_rom <= {16'd7763, 16'd31834};
                15'd2496 : data_rom <= {16'd7766, 16'd31834};
                15'd2497 : data_rom <= {16'd7769, 16'd31833};
                15'd2498 : data_rom <= {16'd7772, 16'd31832};
                15'd2499 : data_rom <= {16'd7775, 16'd31832};
                15'd2500 : data_rom <= {16'd7778, 16'd31831};
                15'd2501 : data_rom <= {16'd7782, 16'd31830};
                15'd2502 : data_rom <= {16'd7785, 16'd31829};
                15'd2503 : data_rom <= {16'd7788, 16'd31829};
                15'd2504 : data_rom <= {16'd7791, 16'd31828};
                15'd2505 : data_rom <= {16'd7794, 16'd31827};
                15'd2506 : data_rom <= {16'd7797, 16'd31826};
                15'd2507 : data_rom <= {16'd7800, 16'd31826};
                15'd2508 : data_rom <= {16'd7803, 16'd31825};
                15'd2509 : data_rom <= {16'd7806, 16'd31824};
                15'd2510 : data_rom <= {16'd7809, 16'd31823};
                15'd2511 : data_rom <= {16'd7812, 16'd31823};
                15'd2512 : data_rom <= {16'd7815, 16'd31822};
                15'd2513 : data_rom <= {16'd7818, 16'd31821};
                15'd2514 : data_rom <= {16'd7821, 16'd31820};
                15'd2515 : data_rom <= {16'd7824, 16'd31820};
                15'd2516 : data_rom <= {16'd7827, 16'd31819};
                15'd2517 : data_rom <= {16'd7830, 16'd31818};
                15'd2518 : data_rom <= {16'd7833, 16'd31817};
                15'd2519 : data_rom <= {16'd7836, 16'd31817};
                15'd2520 : data_rom <= {16'd7840, 16'd31816};
                15'd2521 : data_rom <= {16'd7843, 16'd31815};
                15'd2522 : data_rom <= {16'd7846, 16'd31814};
                15'd2523 : data_rom <= {16'd7849, 16'd31814};
                15'd2524 : data_rom <= {16'd7852, 16'd31813};
                15'd2525 : data_rom <= {16'd7855, 16'd31812};
                15'd2526 : data_rom <= {16'd7858, 16'd31811};
                15'd2527 : data_rom <= {16'd7861, 16'd31811};
                15'd2528 : data_rom <= {16'd7864, 16'd31810};
                15'd2529 : data_rom <= {16'd7867, 16'd31809};
                15'd2530 : data_rom <= {16'd7870, 16'd31808};
                15'd2531 : data_rom <= {16'd7873, 16'd31808};
                15'd2532 : data_rom <= {16'd7876, 16'd31807};
                15'd2533 : data_rom <= {16'd7879, 16'd31806};
                15'd2534 : data_rom <= {16'd7882, 16'd31805};
                15'd2535 : data_rom <= {16'd7885, 16'd31804};
                15'd2536 : data_rom <= {16'd7888, 16'd31804};
                15'd2537 : data_rom <= {16'd7891, 16'd31803};
                15'd2538 : data_rom <= {16'd7894, 16'd31802};
                15'd2539 : data_rom <= {16'd7897, 16'd31801};
                15'd2540 : data_rom <= {16'd7901, 16'd31801};
                15'd2541 : data_rom <= {16'd7904, 16'd31800};
                15'd2542 : data_rom <= {16'd7907, 16'd31799};
                15'd2543 : data_rom <= {16'd7910, 16'd31798};
                15'd2544 : data_rom <= {16'd7913, 16'd31798};
                15'd2545 : data_rom <= {16'd7916, 16'd31797};
                15'd2546 : data_rom <= {16'd7919, 16'd31796};
                15'd2547 : data_rom <= {16'd7922, 16'd31795};
                15'd2548 : data_rom <= {16'd7925, 16'd31795};
                15'd2549 : data_rom <= {16'd7928, 16'd31794};
                15'd2550 : data_rom <= {16'd7931, 16'd31793};
                15'd2551 : data_rom <= {16'd7934, 16'd31792};
                15'd2552 : data_rom <= {16'd7937, 16'd31792};
                15'd2553 : data_rom <= {16'd7940, 16'd31791};
                15'd2554 : data_rom <= {16'd7943, 16'd31790};
                15'd2555 : data_rom <= {16'd7946, 16'd31789};
                15'd2556 : data_rom <= {16'd7949, 16'd31789};
                15'd2557 : data_rom <= {16'd7952, 16'd31788};
                15'd2558 : data_rom <= {16'd7955, 16'd31787};
                15'd2559 : data_rom <= {16'd7958, 16'd31786};
                15'd2560 : data_rom <= {16'd7961, 16'd31785};
                15'd2561 : data_rom <= {16'd7965, 16'd31785};
                15'd2562 : data_rom <= {16'd7968, 16'd31784};
                15'd2563 : data_rom <= {16'd7971, 16'd31783};
                15'd2564 : data_rom <= {16'd7974, 16'd31782};
                15'd2565 : data_rom <= {16'd7977, 16'd31782};
                15'd2566 : data_rom <= {16'd7980, 16'd31781};
                15'd2567 : data_rom <= {16'd7983, 16'd31780};
                15'd2568 : data_rom <= {16'd7986, 16'd31779};
                15'd2569 : data_rom <= {16'd7989, 16'd31779};
                15'd2570 : data_rom <= {16'd7992, 16'd31778};
                15'd2571 : data_rom <= {16'd7995, 16'd31777};
                15'd2572 : data_rom <= {16'd7998, 16'd31776};
                15'd2573 : data_rom <= {16'd8001, 16'd31776};
                15'd2574 : data_rom <= {16'd8004, 16'd31775};
                15'd2575 : data_rom <= {16'd8007, 16'd31774};
                15'd2576 : data_rom <= {16'd8010, 16'd31773};
                15'd2577 : data_rom <= {16'd8013, 16'd31772};
                15'd2578 : data_rom <= {16'd8016, 16'd31772};
                15'd2579 : data_rom <= {16'd8019, 16'd31771};
                15'd2580 : data_rom <= {16'd8022, 16'd31770};
                15'd2581 : data_rom <= {16'd8025, 16'd31769};
                15'd2582 : data_rom <= {16'd8028, 16'd31769};
                15'd2583 : data_rom <= {16'd8032, 16'd31768};
                15'd2584 : data_rom <= {16'd8035, 16'd31767};
                15'd2585 : data_rom <= {16'd8038, 16'd31766};
                15'd2586 : data_rom <= {16'd8041, 16'd31766};
                15'd2587 : data_rom <= {16'd8044, 16'd31765};
                15'd2588 : data_rom <= {16'd8047, 16'd31764};
                15'd2589 : data_rom <= {16'd8050, 16'd31763};
                15'd2590 : data_rom <= {16'd8053, 16'd31762};
                15'd2591 : data_rom <= {16'd8056, 16'd31762};
                15'd2592 : data_rom <= {16'd8059, 16'd31761};
                15'd2593 : data_rom <= {16'd8062, 16'd31760};
                15'd2594 : data_rom <= {16'd8065, 16'd31759};
                15'd2595 : data_rom <= {16'd8068, 16'd31759};
                15'd2596 : data_rom <= {16'd8071, 16'd31758};
                15'd2597 : data_rom <= {16'd8074, 16'd31757};
                15'd2598 : data_rom <= {16'd8077, 16'd31756};
                15'd2599 : data_rom <= {16'd8080, 16'd31755};
                15'd2600 : data_rom <= {16'd8083, 16'd31755};
                15'd2601 : data_rom <= {16'd8086, 16'd31754};
                15'd2602 : data_rom <= {16'd8089, 16'd31753};
                15'd2603 : data_rom <= {16'd8092, 16'd31752};
                15'd2604 : data_rom <= {16'd8095, 16'd31752};
                15'd2605 : data_rom <= {16'd8099, 16'd31751};
                15'd2606 : data_rom <= {16'd8102, 16'd31750};
                15'd2607 : data_rom <= {16'd8105, 16'd31749};
                15'd2608 : data_rom <= {16'd8108, 16'd31749};
                15'd2609 : data_rom <= {16'd8111, 16'd31748};
                15'd2610 : data_rom <= {16'd8114, 16'd31747};
                15'd2611 : data_rom <= {16'd8117, 16'd31746};
                15'd2612 : data_rom <= {16'd8120, 16'd31745};
                15'd2613 : data_rom <= {16'd8123, 16'd31745};
                15'd2614 : data_rom <= {16'd8126, 16'd31744};
                15'd2615 : data_rom <= {16'd8129, 16'd31743};
                15'd2616 : data_rom <= {16'd8132, 16'd31742};
                15'd2617 : data_rom <= {16'd8135, 16'd31742};
                15'd2618 : data_rom <= {16'd8138, 16'd31741};
                15'd2619 : data_rom <= {16'd8141, 16'd31740};
                15'd2620 : data_rom <= {16'd8144, 16'd31739};
                15'd2621 : data_rom <= {16'd8147, 16'd31738};
                15'd2622 : data_rom <= {16'd8150, 16'd31738};
                15'd2623 : data_rom <= {16'd8153, 16'd31737};
                15'd2624 : data_rom <= {16'd8156, 16'd31736};
                15'd2625 : data_rom <= {16'd8159, 16'd31735};
                15'd2626 : data_rom <= {16'd8162, 16'd31734};
                15'd2627 : data_rom <= {16'd8165, 16'd31734};
                15'd2628 : data_rom <= {16'd8169, 16'd31733};
                15'd2629 : data_rom <= {16'd8172, 16'd31732};
                15'd2630 : data_rom <= {16'd8175, 16'd31731};
                15'd2631 : data_rom <= {16'd8178, 16'd31731};
                15'd2632 : data_rom <= {16'd8181, 16'd31730};
                15'd2633 : data_rom <= {16'd8184, 16'd31729};
                15'd2634 : data_rom <= {16'd8187, 16'd31728};
                15'd2635 : data_rom <= {16'd8190, 16'd31727};
                15'd2636 : data_rom <= {16'd8193, 16'd31727};
                15'd2637 : data_rom <= {16'd8196, 16'd31726};
                15'd2638 : data_rom <= {16'd8199, 16'd31725};
                15'd2639 : data_rom <= {16'd8202, 16'd31724};
                15'd2640 : data_rom <= {16'd8205, 16'd31723};
                15'd2641 : data_rom <= {16'd8208, 16'd31723};
                15'd2642 : data_rom <= {16'd8211, 16'd31722};
                15'd2643 : data_rom <= {16'd8214, 16'd31721};
                15'd2644 : data_rom <= {16'd8217, 16'd31720};
                15'd2645 : data_rom <= {16'd8220, 16'd31720};
                15'd2646 : data_rom <= {16'd8223, 16'd31719};
                15'd2647 : data_rom <= {16'd8226, 16'd31718};
                15'd2648 : data_rom <= {16'd8229, 16'd31717};
                15'd2649 : data_rom <= {16'd8232, 16'd31716};
                15'd2650 : data_rom <= {16'd8235, 16'd31716};
                15'd2651 : data_rom <= {16'd8238, 16'd31715};
                15'd2652 : data_rom <= {16'd8242, 16'd31714};
                15'd2653 : data_rom <= {16'd8245, 16'd31713};
                15'd2654 : data_rom <= {16'd8248, 16'd31712};
                15'd2655 : data_rom <= {16'd8251, 16'd31712};
                15'd2656 : data_rom <= {16'd8254, 16'd31711};
                15'd2657 : data_rom <= {16'd8257, 16'd31710};
                15'd2658 : data_rom <= {16'd8260, 16'd31709};
                15'd2659 : data_rom <= {16'd8263, 16'd31708};
                15'd2660 : data_rom <= {16'd8266, 16'd31708};
                15'd2661 : data_rom <= {16'd8269, 16'd31707};
                15'd2662 : data_rom <= {16'd8272, 16'd31706};
                15'd2663 : data_rom <= {16'd8275, 16'd31705};
                15'd2664 : data_rom <= {16'd8278, 16'd31705};
                15'd2665 : data_rom <= {16'd8281, 16'd31704};
                15'd2666 : data_rom <= {16'd8284, 16'd31703};
                15'd2667 : data_rom <= {16'd8287, 16'd31702};
                15'd2668 : data_rom <= {16'd8290, 16'd31701};
                15'd2669 : data_rom <= {16'd8293, 16'd31701};
                15'd2670 : data_rom <= {16'd8296, 16'd31700};
                15'd2671 : data_rom <= {16'd8299, 16'd31699};
                15'd2672 : data_rom <= {16'd8302, 16'd31698};
                15'd2673 : data_rom <= {16'd8305, 16'd31697};
                15'd2674 : data_rom <= {16'd8308, 16'd31697};
                15'd2675 : data_rom <= {16'd8311, 16'd31696};
                15'd2676 : data_rom <= {16'd8314, 16'd31695};
                15'd2677 : data_rom <= {16'd8318, 16'd31694};
                15'd2678 : data_rom <= {16'd8321, 16'd31693};
                15'd2679 : data_rom <= {16'd8324, 16'd31693};
                15'd2680 : data_rom <= {16'd8327, 16'd31692};
                15'd2681 : data_rom <= {16'd8330, 16'd31691};
                15'd2682 : data_rom <= {16'd8333, 16'd31690};
                15'd2683 : data_rom <= {16'd8336, 16'd31689};
                15'd2684 : data_rom <= {16'd8339, 16'd31689};
                15'd2685 : data_rom <= {16'd8342, 16'd31688};
                15'd2686 : data_rom <= {16'd8345, 16'd31687};
                15'd2687 : data_rom <= {16'd8348, 16'd31686};
                15'd2688 : data_rom <= {16'd8351, 16'd31685};
                15'd2689 : data_rom <= {16'd8354, 16'd31685};
                15'd2690 : data_rom <= {16'd8357, 16'd31684};
                15'd2691 : data_rom <= {16'd8360, 16'd31683};
                15'd2692 : data_rom <= {16'd8363, 16'd31682};
                15'd2693 : data_rom <= {16'd8366, 16'd31681};
                15'd2694 : data_rom <= {16'd8369, 16'd31681};
                15'd2695 : data_rom <= {16'd8372, 16'd31680};
                15'd2696 : data_rom <= {16'd8375, 16'd31679};
                15'd2697 : data_rom <= {16'd8378, 16'd31678};
                15'd2698 : data_rom <= {16'd8381, 16'd31677};
                15'd2699 : data_rom <= {16'd8384, 16'd31677};
                15'd2700 : data_rom <= {16'd8387, 16'd31676};
                15'd2701 : data_rom <= {16'd8390, 16'd31675};
                15'd2702 : data_rom <= {16'd8393, 16'd31674};
                15'd2703 : data_rom <= {16'd8396, 16'd31673};
                15'd2704 : data_rom <= {16'd8400, 16'd31673};
                15'd2705 : data_rom <= {16'd8403, 16'd31672};
                15'd2706 : data_rom <= {16'd8406, 16'd31671};
                15'd2707 : data_rom <= {16'd8409, 16'd31670};
                15'd2708 : data_rom <= {16'd8412, 16'd31669};
                15'd2709 : data_rom <= {16'd8415, 16'd31669};
                15'd2710 : data_rom <= {16'd8418, 16'd31668};
                15'd2711 : data_rom <= {16'd8421, 16'd31667};
                15'd2712 : data_rom <= {16'd8424, 16'd31666};
                15'd2713 : data_rom <= {16'd8427, 16'd31665};
                15'd2714 : data_rom <= {16'd8430, 16'd31664};
                15'd2715 : data_rom <= {16'd8433, 16'd31664};
                15'd2716 : data_rom <= {16'd8436, 16'd31663};
                15'd2717 : data_rom <= {16'd8439, 16'd31662};
                15'd2718 : data_rom <= {16'd8442, 16'd31661};
                15'd2719 : data_rom <= {16'd8445, 16'd31660};
                15'd2720 : data_rom <= {16'd8448, 16'd31660};
                15'd2721 : data_rom <= {16'd8451, 16'd31659};
                15'd2722 : data_rom <= {16'd8454, 16'd31658};
                15'd2723 : data_rom <= {16'd8457, 16'd31657};
                15'd2724 : data_rom <= {16'd8460, 16'd31656};
                15'd2725 : data_rom <= {16'd8463, 16'd31656};
                15'd2726 : data_rom <= {16'd8466, 16'd31655};
                15'd2727 : data_rom <= {16'd8469, 16'd31654};
                15'd2728 : data_rom <= {16'd8472, 16'd31653};
                15'd2729 : data_rom <= {16'd8475, 16'd31652};
                15'd2730 : data_rom <= {16'd8478, 16'd31652};
                15'd2731 : data_rom <= {16'd8481, 16'd31651};
                15'd2732 : data_rom <= {16'd8485, 16'd31650};
                15'd2733 : data_rom <= {16'd8488, 16'd31649};
                15'd2734 : data_rom <= {16'd8491, 16'd31648};
                15'd2735 : data_rom <= {16'd8494, 16'd31647};
                15'd2736 : data_rom <= {16'd8497, 16'd31647};
                15'd2737 : data_rom <= {16'd8500, 16'd31646};
                15'd2738 : data_rom <= {16'd8503, 16'd31645};
                15'd2739 : data_rom <= {16'd8506, 16'd31644};
                15'd2740 : data_rom <= {16'd8509, 16'd31643};
                15'd2741 : data_rom <= {16'd8512, 16'd31643};
                15'd2742 : data_rom <= {16'd8515, 16'd31642};
                15'd2743 : data_rom <= {16'd8518, 16'd31641};
                15'd2744 : data_rom <= {16'd8521, 16'd31640};
                15'd2745 : data_rom <= {16'd8524, 16'd31639};
                15'd2746 : data_rom <= {16'd8527, 16'd31638};
                15'd2747 : data_rom <= {16'd8530, 16'd31638};
                15'd2748 : data_rom <= {16'd8533, 16'd31637};
                15'd2749 : data_rom <= {16'd8536, 16'd31636};
                15'd2750 : data_rom <= {16'd8539, 16'd31635};
                15'd2751 : data_rom <= {16'd8542, 16'd31634};
                15'd2752 : data_rom <= {16'd8545, 16'd31634};
                15'd2753 : data_rom <= {16'd8548, 16'd31633};
                15'd2754 : data_rom <= {16'd8551, 16'd31632};
                15'd2755 : data_rom <= {16'd8554, 16'd31631};
                15'd2756 : data_rom <= {16'd8557, 16'd31630};
                15'd2757 : data_rom <= {16'd8560, 16'd31629};
                15'd2758 : data_rom <= {16'd8563, 16'd31629};
                15'd2759 : data_rom <= {16'd8566, 16'd31628};
                15'd2760 : data_rom <= {16'd8569, 16'd31627};
                15'd2761 : data_rom <= {16'd8572, 16'd31626};
                15'd2762 : data_rom <= {16'd8576, 16'd31625};
                15'd2763 : data_rom <= {16'd8579, 16'd31625};
                15'd2764 : data_rom <= {16'd8582, 16'd31624};
                15'd2765 : data_rom <= {16'd8585, 16'd31623};
                15'd2766 : data_rom <= {16'd8588, 16'd31622};
                15'd2767 : data_rom <= {16'd8591, 16'd31621};
                15'd2768 : data_rom <= {16'd8594, 16'd31620};
                15'd2769 : data_rom <= {16'd8597, 16'd31620};
                15'd2770 : data_rom <= {16'd8600, 16'd31619};
                15'd2771 : data_rom <= {16'd8603, 16'd31618};
                15'd2772 : data_rom <= {16'd8606, 16'd31617};
                15'd2773 : data_rom <= {16'd8609, 16'd31616};
                15'd2774 : data_rom <= {16'd8612, 16'd31615};
                15'd2775 : data_rom <= {16'd8615, 16'd31615};
                15'd2776 : data_rom <= {16'd8618, 16'd31614};
                15'd2777 : data_rom <= {16'd8621, 16'd31613};
                15'd2778 : data_rom <= {16'd8624, 16'd31612};
                15'd2779 : data_rom <= {16'd8627, 16'd31611};
                15'd2780 : data_rom <= {16'd8630, 16'd31610};
                15'd2781 : data_rom <= {16'd8633, 16'd31610};
                15'd2782 : data_rom <= {16'd8636, 16'd31609};
                15'd2783 : data_rom <= {16'd8639, 16'd31608};
                15'd2784 : data_rom <= {16'd8642, 16'd31607};
                15'd2785 : data_rom <= {16'd8645, 16'd31606};
                15'd2786 : data_rom <= {16'd8648, 16'd31606};
                15'd2787 : data_rom <= {16'd8651, 16'd31605};
                15'd2788 : data_rom <= {16'd8654, 16'd31604};
                15'd2789 : data_rom <= {16'd8657, 16'd31603};
                15'd2790 : data_rom <= {16'd8660, 16'd31602};
                15'd2791 : data_rom <= {16'd8663, 16'd31601};
                15'd2792 : data_rom <= {16'd8666, 16'd31601};
                15'd2793 : data_rom <= {16'd8669, 16'd31600};
                15'd2794 : data_rom <= {16'd8673, 16'd31599};
                15'd2795 : data_rom <= {16'd8676, 16'd31598};
                15'd2796 : data_rom <= {16'd8679, 16'd31597};
                15'd2797 : data_rom <= {16'd8682, 16'd31596};
                15'd2798 : data_rom <= {16'd8685, 16'd31596};
                15'd2799 : data_rom <= {16'd8688, 16'd31595};
                15'd2800 : data_rom <= {16'd8691, 16'd31594};
                15'd2801 : data_rom <= {16'd8694, 16'd31593};
                15'd2802 : data_rom <= {16'd8697, 16'd31592};
                15'd2803 : data_rom <= {16'd8700, 16'd31591};
                15'd2804 : data_rom <= {16'd8703, 16'd31591};
                15'd2805 : data_rom <= {16'd8706, 16'd31590};
                15'd2806 : data_rom <= {16'd8709, 16'd31589};
                15'd2807 : data_rom <= {16'd8712, 16'd31588};
                15'd2808 : data_rom <= {16'd8715, 16'd31587};
                15'd2809 : data_rom <= {16'd8718, 16'd31586};
                15'd2810 : data_rom <= {16'd8721, 16'd31586};
                15'd2811 : data_rom <= {16'd8724, 16'd31585};
                15'd2812 : data_rom <= {16'd8727, 16'd31584};
                15'd2813 : data_rom <= {16'd8730, 16'd31583};
                15'd2814 : data_rom <= {16'd8733, 16'd31582};
                15'd2815 : data_rom <= {16'd8736, 16'd31581};
                15'd2816 : data_rom <= {16'd8739, 16'd31581};
                15'd2817 : data_rom <= {16'd8742, 16'd31580};
                15'd2818 : data_rom <= {16'd8745, 16'd31579};
                15'd2819 : data_rom <= {16'd8748, 16'd31578};
                15'd2820 : data_rom <= {16'd8751, 16'd31577};
                15'd2821 : data_rom <= {16'd8754, 16'd31576};
                15'd2822 : data_rom <= {16'd8757, 16'd31575};
                15'd2823 : data_rom <= {16'd8760, 16'd31575};
                15'd2824 : data_rom <= {16'd8763, 16'd31574};
                15'd2825 : data_rom <= {16'd8766, 16'd31573};
                15'd2826 : data_rom <= {16'd8769, 16'd31572};
                15'd2827 : data_rom <= {16'd8772, 16'd31571};
                15'd2828 : data_rom <= {16'd8775, 16'd31570};
                15'd2829 : data_rom <= {16'd8778, 16'd31570};
                15'd2830 : data_rom <= {16'd8782, 16'd31569};
                15'd2831 : data_rom <= {16'd8785, 16'd31568};
                15'd2832 : data_rom <= {16'd8788, 16'd31567};
                15'd2833 : data_rom <= {16'd8791, 16'd31566};
                15'd2834 : data_rom <= {16'd8794, 16'd31565};
                15'd2835 : data_rom <= {16'd8797, 16'd31565};
                15'd2836 : data_rom <= {16'd8800, 16'd31564};
                15'd2837 : data_rom <= {16'd8803, 16'd31563};
                15'd2838 : data_rom <= {16'd8806, 16'd31562};
                15'd2839 : data_rom <= {16'd8809, 16'd31561};
                15'd2840 : data_rom <= {16'd8812, 16'd31560};
                15'd2841 : data_rom <= {16'd8815, 16'd31559};
                15'd2842 : data_rom <= {16'd8818, 16'd31559};
                15'd2843 : data_rom <= {16'd8821, 16'd31558};
                15'd2844 : data_rom <= {16'd8824, 16'd31557};
                15'd2845 : data_rom <= {16'd8827, 16'd31556};
                15'd2846 : data_rom <= {16'd8830, 16'd31555};
                15'd2847 : data_rom <= {16'd8833, 16'd31554};
                15'd2848 : data_rom <= {16'd8836, 16'd31554};
                15'd2849 : data_rom <= {16'd8839, 16'd31553};
                15'd2850 : data_rom <= {16'd8842, 16'd31552};
                15'd2851 : data_rom <= {16'd8845, 16'd31551};
                15'd2852 : data_rom <= {16'd8848, 16'd31550};
                15'd2853 : data_rom <= {16'd8851, 16'd31549};
                15'd2854 : data_rom <= {16'd8854, 16'd31548};
                15'd2855 : data_rom <= {16'd8857, 16'd31548};
                15'd2856 : data_rom <= {16'd8860, 16'd31547};
                15'd2857 : data_rom <= {16'd8863, 16'd31546};
                15'd2858 : data_rom <= {16'd8866, 16'd31545};
                15'd2859 : data_rom <= {16'd8869, 16'd31544};
                15'd2860 : data_rom <= {16'd8872, 16'd31543};
                15'd2861 : data_rom <= {16'd8875, 16'd31543};
                15'd2862 : data_rom <= {16'd8878, 16'd31542};
                15'd2863 : data_rom <= {16'd8881, 16'd31541};
                15'd2864 : data_rom <= {16'd8884, 16'd31540};
                15'd2865 : data_rom <= {16'd8887, 16'd31539};
                15'd2866 : data_rom <= {16'd8890, 16'd31538};
                15'd2867 : data_rom <= {16'd8893, 16'd31537};
                15'd2868 : data_rom <= {16'd8896, 16'd31537};
                15'd2869 : data_rom <= {16'd8899, 16'd31536};
                15'd2870 : data_rom <= {16'd8903, 16'd31535};
                15'd2871 : data_rom <= {16'd8906, 16'd31534};
                15'd2872 : data_rom <= {16'd8909, 16'd31533};
                15'd2873 : data_rom <= {16'd8912, 16'd31532};
                15'd2874 : data_rom <= {16'd8915, 16'd31531};
                15'd2875 : data_rom <= {16'd8918, 16'd31531};
                15'd2876 : data_rom <= {16'd8921, 16'd31530};
                15'd2877 : data_rom <= {16'd8924, 16'd31529};
                15'd2878 : data_rom <= {16'd8927, 16'd31528};
                15'd2879 : data_rom <= {16'd8930, 16'd31527};
                15'd2880 : data_rom <= {16'd8933, 16'd31526};
                15'd2881 : data_rom <= {16'd8936, 16'd31525};
                15'd2882 : data_rom <= {16'd8939, 16'd31525};
                15'd2883 : data_rom <= {16'd8942, 16'd31524};
                15'd2884 : data_rom <= {16'd8945, 16'd31523};
                15'd2885 : data_rom <= {16'd8948, 16'd31522};
                15'd2886 : data_rom <= {16'd8951, 16'd31521};
                15'd2887 : data_rom <= {16'd8954, 16'd31520};
                15'd2888 : data_rom <= {16'd8957, 16'd31519};
                15'd2889 : data_rom <= {16'd8960, 16'd31519};
                15'd2890 : data_rom <= {16'd8963, 16'd31518};
                15'd2891 : data_rom <= {16'd8966, 16'd31517};
                15'd2892 : data_rom <= {16'd8969, 16'd31516};
                15'd2893 : data_rom <= {16'd8972, 16'd31515};
                15'd2894 : data_rom <= {16'd8975, 16'd31514};
                15'd2895 : data_rom <= {16'd8978, 16'd31513};
                15'd2896 : data_rom <= {16'd8981, 16'd31513};
                15'd2897 : data_rom <= {16'd8984, 16'd31512};
                15'd2898 : data_rom <= {16'd8987, 16'd31511};
                15'd2899 : data_rom <= {16'd8990, 16'd31510};
                15'd2900 : data_rom <= {16'd8993, 16'd31509};
                15'd2901 : data_rom <= {16'd8996, 16'd31508};
                15'd2902 : data_rom <= {16'd8999, 16'd31507};
                15'd2903 : data_rom <= {16'd9002, 16'd31507};
                15'd2904 : data_rom <= {16'd9005, 16'd31506};
                15'd2905 : data_rom <= {16'd9008, 16'd31505};
                15'd2906 : data_rom <= {16'd9011, 16'd31504};
                15'd2907 : data_rom <= {16'd9014, 16'd31503};
                15'd2908 : data_rom <= {16'd9017, 16'd31502};
                15'd2909 : data_rom <= {16'd9020, 16'd31501};
                15'd2910 : data_rom <= {16'd9023, 16'd31500};
                15'd2911 : data_rom <= {16'd9026, 16'd31500};
                15'd2912 : data_rom <= {16'd9029, 16'd31499};
                15'd2913 : data_rom <= {16'd9032, 16'd31498};
                15'd2914 : data_rom <= {16'd9035, 16'd31497};
                15'd2915 : data_rom <= {16'd9038, 16'd31496};
                15'd2916 : data_rom <= {16'd9042, 16'd31495};
                15'd2917 : data_rom <= {16'd9045, 16'd31494};
                15'd2918 : data_rom <= {16'd9048, 16'd31494};
                15'd2919 : data_rom <= {16'd9051, 16'd31493};
                15'd2920 : data_rom <= {16'd9054, 16'd31492};
                15'd2921 : data_rom <= {16'd9057, 16'd31491};
                15'd2922 : data_rom <= {16'd9060, 16'd31490};
                15'd2923 : data_rom <= {16'd9063, 16'd31489};
                15'd2924 : data_rom <= {16'd9066, 16'd31488};
                15'd2925 : data_rom <= {16'd9069, 16'd31487};
                15'd2926 : data_rom <= {16'd9072, 16'd31487};
                15'd2927 : data_rom <= {16'd9075, 16'd31486};
                15'd2928 : data_rom <= {16'd9078, 16'd31485};
                15'd2929 : data_rom <= {16'd9081, 16'd31484};
                15'd2930 : data_rom <= {16'd9084, 16'd31483};
                15'd2931 : data_rom <= {16'd9087, 16'd31482};
                15'd2932 : data_rom <= {16'd9090, 16'd31481};
                15'd2933 : data_rom <= {16'd9093, 16'd31480};
                15'd2934 : data_rom <= {16'd9096, 16'd31480};
                15'd2935 : data_rom <= {16'd9099, 16'd31479};
                15'd2936 : data_rom <= {16'd9102, 16'd31478};
                15'd2937 : data_rom <= {16'd9105, 16'd31477};
                15'd2938 : data_rom <= {16'd9108, 16'd31476};
                15'd2939 : data_rom <= {16'd9111, 16'd31475};
                15'd2940 : data_rom <= {16'd9114, 16'd31474};
                15'd2941 : data_rom <= {16'd9117, 16'd31474};
                15'd2942 : data_rom <= {16'd9120, 16'd31473};
                15'd2943 : data_rom <= {16'd9123, 16'd31472};
                15'd2944 : data_rom <= {16'd9126, 16'd31471};
                15'd2945 : data_rom <= {16'd9129, 16'd31470};
                15'd2946 : data_rom <= {16'd9132, 16'd31469};
                15'd2947 : data_rom <= {16'd9135, 16'd31468};
                15'd2948 : data_rom <= {16'd9138, 16'd31467};
                15'd2949 : data_rom <= {16'd9141, 16'd31467};
                15'd2950 : data_rom <= {16'd9144, 16'd31466};
                15'd2951 : data_rom <= {16'd9147, 16'd31465};
                15'd2952 : data_rom <= {16'd9150, 16'd31464};
                15'd2953 : data_rom <= {16'd9153, 16'd31463};
                15'd2954 : data_rom <= {16'd9156, 16'd31462};
                15'd2955 : data_rom <= {16'd9159, 16'd31461};
                15'd2956 : data_rom <= {16'd9162, 16'd31460};
                15'd2957 : data_rom <= {16'd9165, 16'd31459};
                15'd2958 : data_rom <= {16'd9168, 16'd31459};
                15'd2959 : data_rom <= {16'd9171, 16'd31458};
                15'd2960 : data_rom <= {16'd9174, 16'd31457};
                15'd2961 : data_rom <= {16'd9177, 16'd31456};
                15'd2962 : data_rom <= {16'd9180, 16'd31455};
                15'd2963 : data_rom <= {16'd9183, 16'd31454};
                15'd2964 : data_rom <= {16'd9186, 16'd31453};
                15'd2965 : data_rom <= {16'd9189, 16'd31452};
                15'd2966 : data_rom <= {16'd9192, 16'd31452};
                15'd2967 : data_rom <= {16'd9195, 16'd31451};
                15'd2968 : data_rom <= {16'd9198, 16'd31450};
                15'd2969 : data_rom <= {16'd9201, 16'd31449};
                15'd2970 : data_rom <= {16'd9204, 16'd31448};
                15'd2971 : data_rom <= {16'd9207, 16'd31447};
                15'd2972 : data_rom <= {16'd9210, 16'd31446};
                15'd2973 : data_rom <= {16'd9213, 16'd31445};
                15'd2974 : data_rom <= {16'd9217, 16'd31445};
                15'd2975 : data_rom <= {16'd9220, 16'd31444};
                15'd2976 : data_rom <= {16'd9223, 16'd31443};
                15'd2977 : data_rom <= {16'd9226, 16'd31442};
                15'd2978 : data_rom <= {16'd9229, 16'd31441};
                15'd2979 : data_rom <= {16'd9232, 16'd31440};
                15'd2980 : data_rom <= {16'd9235, 16'd31439};
                15'd2981 : data_rom <= {16'd9238, 16'd31438};
                15'd2982 : data_rom <= {16'd9241, 16'd31437};
                15'd2983 : data_rom <= {16'd9244, 16'd31437};
                15'd2984 : data_rom <= {16'd9247, 16'd31436};
                15'd2985 : data_rom <= {16'd9250, 16'd31435};
                15'd2986 : data_rom <= {16'd9253, 16'd31434};
                15'd2987 : data_rom <= {16'd9256, 16'd31433};
                15'd2988 : data_rom <= {16'd9259, 16'd31432};
                15'd2989 : data_rom <= {16'd9262, 16'd31431};
                15'd2990 : data_rom <= {16'd9265, 16'd31430};
                15'd2991 : data_rom <= {16'd9268, 16'd31429};
                15'd2992 : data_rom <= {16'd9271, 16'd31429};
                15'd2993 : data_rom <= {16'd9274, 16'd31428};
                15'd2994 : data_rom <= {16'd9277, 16'd31427};
                15'd2995 : data_rom <= {16'd9280, 16'd31426};
                15'd2996 : data_rom <= {16'd9283, 16'd31425};
                15'd2997 : data_rom <= {16'd9286, 16'd31424};
                15'd2998 : data_rom <= {16'd9289, 16'd31423};
                15'd2999 : data_rom <= {16'd9292, 16'd31422};
                15'd3000 : data_rom <= {16'd9295, 16'd31421};
                15'd3001 : data_rom <= {16'd9298, 16'd31421};
                15'd3002 : data_rom <= {16'd9301, 16'd31420};
                15'd3003 : data_rom <= {16'd9304, 16'd31419};
                15'd3004 : data_rom <= {16'd9307, 16'd31418};
                15'd3005 : data_rom <= {16'd9310, 16'd31417};
                15'd3006 : data_rom <= {16'd9313, 16'd31416};
                15'd3007 : data_rom <= {16'd9316, 16'd31415};
                15'd3008 : data_rom <= {16'd9319, 16'd31414};
                15'd3009 : data_rom <= {16'd9322, 16'd31413};
                15'd3010 : data_rom <= {16'd9325, 16'd31413};
                15'd3011 : data_rom <= {16'd9328, 16'd31412};
                15'd3012 : data_rom <= {16'd9331, 16'd31411};
                15'd3013 : data_rom <= {16'd9334, 16'd31410};
                15'd3014 : data_rom <= {16'd9337, 16'd31409};
                15'd3015 : data_rom <= {16'd9340, 16'd31408};
                15'd3016 : data_rom <= {16'd9343, 16'd31407};
                15'd3017 : data_rom <= {16'd9346, 16'd31406};
                15'd3018 : data_rom <= {16'd9349, 16'd31405};
                15'd3019 : data_rom <= {16'd9352, 16'd31404};
                15'd3020 : data_rom <= {16'd9355, 16'd31404};
                15'd3021 : data_rom <= {16'd9358, 16'd31403};
                15'd3022 : data_rom <= {16'd9361, 16'd31402};
                15'd3023 : data_rom <= {16'd9364, 16'd31401};
                15'd3024 : data_rom <= {16'd9367, 16'd31400};
                15'd3025 : data_rom <= {16'd9370, 16'd31399};
                15'd3026 : data_rom <= {16'd9373, 16'd31398};
                15'd3027 : data_rom <= {16'd9376, 16'd31397};
                15'd3028 : data_rom <= {16'd9379, 16'd31396};
                15'd3029 : data_rom <= {16'd9382, 16'd31395};
                15'd3030 : data_rom <= {16'd9385, 16'd31395};
                15'd3031 : data_rom <= {16'd9388, 16'd31394};
                15'd3032 : data_rom <= {16'd9391, 16'd31393};
                15'd3033 : data_rom <= {16'd9394, 16'd31392};
                15'd3034 : data_rom <= {16'd9397, 16'd31391};
                15'd3035 : data_rom <= {16'd9400, 16'd31390};
                15'd3036 : data_rom <= {16'd9403, 16'd31389};
                15'd3037 : data_rom <= {16'd9406, 16'd31388};
                15'd3038 : data_rom <= {16'd9409, 16'd31387};
                15'd3039 : data_rom <= {16'd9412, 16'd31386};
                15'd3040 : data_rom <= {16'd9415, 16'd31386};
                15'd3041 : data_rom <= {16'd9418, 16'd31385};
                15'd3042 : data_rom <= {16'd9421, 16'd31384};
                15'd3043 : data_rom <= {16'd9424, 16'd31383};
                15'd3044 : data_rom <= {16'd9427, 16'd31382};
                15'd3045 : data_rom <= {16'd9430, 16'd31381};
                15'd3046 : data_rom <= {16'd9433, 16'd31380};
                15'd3047 : data_rom <= {16'd9436, 16'd31379};
                15'd3048 : data_rom <= {16'd9439, 16'd31378};
                15'd3049 : data_rom <= {16'd9442, 16'd31377};
                15'd3050 : data_rom <= {16'd9445, 16'd31377};
                15'd3051 : data_rom <= {16'd9448, 16'd31376};
                15'd3052 : data_rom <= {16'd9451, 16'd31375};
                15'd3053 : data_rom <= {16'd9454, 16'd31374};
                15'd3054 : data_rom <= {16'd9457, 16'd31373};
                15'd3055 : data_rom <= {16'd9460, 16'd31372};
                15'd3056 : data_rom <= {16'd9463, 16'd31371};
                15'd3057 : data_rom <= {16'd9466, 16'd31370};
                15'd3058 : data_rom <= {16'd9469, 16'd31369};
                15'd3059 : data_rom <= {16'd9472, 16'd31368};
                15'd3060 : data_rom <= {16'd9475, 16'd31367};
                15'd3061 : data_rom <= {16'd9478, 16'd31367};
                15'd3062 : data_rom <= {16'd9481, 16'd31366};
                15'd3063 : data_rom <= {16'd9484, 16'd31365};
                15'd3064 : data_rom <= {16'd9487, 16'd31364};
                15'd3065 : data_rom <= {16'd9490, 16'd31363};
                15'd3066 : data_rom <= {16'd9494, 16'd31362};
                15'd3067 : data_rom <= {16'd9497, 16'd31361};
                15'd3068 : data_rom <= {16'd9500, 16'd31360};
                15'd3069 : data_rom <= {16'd9503, 16'd31359};
                15'd3070 : data_rom <= {16'd9506, 16'd31358};
                15'd3071 : data_rom <= {16'd9509, 16'd31357};
                15'd3072 : data_rom <= {16'd9512, 16'd31357};
                15'd3073 : data_rom <= {16'd9515, 16'd31356};
                15'd3074 : data_rom <= {16'd9518, 16'd31355};
                15'd3075 : data_rom <= {16'd9521, 16'd31354};
                15'd3076 : data_rom <= {16'd9524, 16'd31353};
                15'd3077 : data_rom <= {16'd9527, 16'd31352};
                15'd3078 : data_rom <= {16'd9530, 16'd31351};
                15'd3079 : data_rom <= {16'd9533, 16'd31350};
                15'd3080 : data_rom <= {16'd9536, 16'd31349};
                15'd3081 : data_rom <= {16'd9539, 16'd31348};
                15'd3082 : data_rom <= {16'd9542, 16'd31347};
                15'd3083 : data_rom <= {16'd9545, 16'd31346};
                15'd3084 : data_rom <= {16'd9548, 16'd31346};
                15'd3085 : data_rom <= {16'd9551, 16'd31345};
                15'd3086 : data_rom <= {16'd9554, 16'd31344};
                15'd3087 : data_rom <= {16'd9557, 16'd31343};
                15'd3088 : data_rom <= {16'd9560, 16'd31342};
                15'd3089 : data_rom <= {16'd9563, 16'd31341};
                15'd3090 : data_rom <= {16'd9566, 16'd31340};
                15'd3091 : data_rom <= {16'd9569, 16'd31339};
                15'd3092 : data_rom <= {16'd9572, 16'd31338};
                15'd3093 : data_rom <= {16'd9575, 16'd31337};
                15'd3094 : data_rom <= {16'd9578, 16'd31336};
                15'd3095 : data_rom <= {16'd9581, 16'd31335};
                15'd3096 : data_rom <= {16'd9584, 16'd31335};
                15'd3097 : data_rom <= {16'd9587, 16'd31334};
                15'd3098 : data_rom <= {16'd9590, 16'd31333};
                15'd3099 : data_rom <= {16'd9593, 16'd31332};
                15'd3100 : data_rom <= {16'd9596, 16'd31331};
                15'd3101 : data_rom <= {16'd9599, 16'd31330};
                15'd3102 : data_rom <= {16'd9602, 16'd31329};
                15'd3103 : data_rom <= {16'd9605, 16'd31328};
                15'd3104 : data_rom <= {16'd9608, 16'd31327};
                15'd3105 : data_rom <= {16'd9611, 16'd31326};
                15'd3106 : data_rom <= {16'd9614, 16'd31325};
                15'd3107 : data_rom <= {16'd9617, 16'd31324};
                15'd3108 : data_rom <= {16'd9620, 16'd31324};
                15'd3109 : data_rom <= {16'd9623, 16'd31323};
                15'd3110 : data_rom <= {16'd9626, 16'd31322};
                15'd3111 : data_rom <= {16'd9629, 16'd31321};
                15'd3112 : data_rom <= {16'd9632, 16'd31320};
                15'd3113 : data_rom <= {16'd9635, 16'd31319};
                15'd3114 : data_rom <= {16'd9638, 16'd31318};
                15'd3115 : data_rom <= {16'd9641, 16'd31317};
                15'd3116 : data_rom <= {16'd9644, 16'd31316};
                15'd3117 : data_rom <= {16'd9647, 16'd31315};
                15'd3118 : data_rom <= {16'd9650, 16'd31314};
                15'd3119 : data_rom <= {16'd9653, 16'd31313};
                15'd3120 : data_rom <= {16'd9656, 16'd31312};
                15'd3121 : data_rom <= {16'd9659, 16'd31311};
                15'd3122 : data_rom <= {16'd9662, 16'd31311};
                15'd3123 : data_rom <= {16'd9665, 16'd31310};
                15'd3124 : data_rom <= {16'd9668, 16'd31309};
                15'd3125 : data_rom <= {16'd9671, 16'd31308};
                15'd3126 : data_rom <= {16'd9674, 16'd31307};
                15'd3127 : data_rom <= {16'd9677, 16'd31306};
                15'd3128 : data_rom <= {16'd9680, 16'd31305};
                15'd3129 : data_rom <= {16'd9683, 16'd31304};
                15'd3130 : data_rom <= {16'd9686, 16'd31303};
                15'd3131 : data_rom <= {16'd9689, 16'd31302};
                15'd3132 : data_rom <= {16'd9692, 16'd31301};
                15'd3133 : data_rom <= {16'd9695, 16'd31300};
                15'd3134 : data_rom <= {16'd9698, 16'd31299};
                15'd3135 : data_rom <= {16'd9701, 16'd31298};
                15'd3136 : data_rom <= {16'd9704, 16'd31298};
                15'd3137 : data_rom <= {16'd9707, 16'd31297};
                15'd3138 : data_rom <= {16'd9710, 16'd31296};
                15'd3139 : data_rom <= {16'd9713, 16'd31295};
                15'd3140 : data_rom <= {16'd9716, 16'd31294};
                15'd3141 : data_rom <= {16'd9719, 16'd31293};
                15'd3142 : data_rom <= {16'd9722, 16'd31292};
                15'd3143 : data_rom <= {16'd9725, 16'd31291};
                15'd3144 : data_rom <= {16'd9728, 16'd31290};
                15'd3145 : data_rom <= {16'd9731, 16'd31289};
                15'd3146 : data_rom <= {16'd9734, 16'd31288};
                15'd3147 : data_rom <= {16'd9737, 16'd31287};
                15'd3148 : data_rom <= {16'd9740, 16'd31286};
                15'd3149 : data_rom <= {16'd9743, 16'd31285};
                15'd3150 : data_rom <= {16'd9746, 16'd31285};
                15'd3151 : data_rom <= {16'd9749, 16'd31284};
                15'd3152 : data_rom <= {16'd9752, 16'd31283};
                15'd3153 : data_rom <= {16'd9755, 16'd31282};
                15'd3154 : data_rom <= {16'd9758, 16'd31281};
                15'd3155 : data_rom <= {16'd9761, 16'd31280};
                15'd3156 : data_rom <= {16'd9764, 16'd31279};
                15'd3157 : data_rom <= {16'd9767, 16'd31278};
                15'd3158 : data_rom <= {16'd9770, 16'd31277};
                15'd3159 : data_rom <= {16'd9773, 16'd31276};
                15'd3160 : data_rom <= {16'd9776, 16'd31275};
                15'd3161 : data_rom <= {16'd9779, 16'd31274};
                15'd3162 : data_rom <= {16'd9782, 16'd31273};
                15'd3163 : data_rom <= {16'd9785, 16'd31272};
                15'd3164 : data_rom <= {16'd9788, 16'd31271};
                15'd3165 : data_rom <= {16'd9791, 16'd31270};
                15'd3166 : data_rom <= {16'd9794, 16'd31270};
                15'd3167 : data_rom <= {16'd9797, 16'd31269};
                15'd3168 : data_rom <= {16'd9800, 16'd31268};
                15'd3169 : data_rom <= {16'd9803, 16'd31267};
                15'd3170 : data_rom <= {16'd9806, 16'd31266};
                15'd3171 : data_rom <= {16'd9809, 16'd31265};
                15'd3172 : data_rom <= {16'd9812, 16'd31264};
                15'd3173 : data_rom <= {16'd9815, 16'd31263};
                15'd3174 : data_rom <= {16'd9818, 16'd31262};
                15'd3175 : data_rom <= {16'd9821, 16'd31261};
                15'd3176 : data_rom <= {16'd9824, 16'd31260};
                15'd3177 : data_rom <= {16'd9827, 16'd31259};
                15'd3178 : data_rom <= {16'd9830, 16'd31258};
                15'd3179 : data_rom <= {16'd9833, 16'd31257};
                15'd3180 : data_rom <= {16'd9836, 16'd31256};
                15'd3181 : data_rom <= {16'd9839, 16'd31255};
                15'd3182 : data_rom <= {16'd9842, 16'd31254};
                15'd3183 : data_rom <= {16'd9845, 16'd31254};
                15'd3184 : data_rom <= {16'd9848, 16'd31253};
                15'd3185 : data_rom <= {16'd9851, 16'd31252};
                15'd3186 : data_rom <= {16'd9854, 16'd31251};
                15'd3187 : data_rom <= {16'd9857, 16'd31250};
                15'd3188 : data_rom <= {16'd9860, 16'd31249};
                15'd3189 : data_rom <= {16'd9863, 16'd31248};
                15'd3190 : data_rom <= {16'd9866, 16'd31247};
                15'd3191 : data_rom <= {16'd9869, 16'd31246};
                15'd3192 : data_rom <= {16'd9872, 16'd31245};
                15'd3193 : data_rom <= {16'd9875, 16'd31244};
                15'd3194 : data_rom <= {16'd9878, 16'd31243};
                15'd3195 : data_rom <= {16'd9881, 16'd31242};
                15'd3196 : data_rom <= {16'd9884, 16'd31241};
                15'd3197 : data_rom <= {16'd9887, 16'd31240};
                15'd3198 : data_rom <= {16'd9890, 16'd31239};
                15'd3199 : data_rom <= {16'd9893, 16'd31238};
                15'd3200 : data_rom <= {16'd9896, 16'd31237};
                15'd3201 : data_rom <= {16'd9899, 16'd31236};
                15'd3202 : data_rom <= {16'd9902, 16'd31236};
                15'd3203 : data_rom <= {16'd9905, 16'd31235};
                15'd3204 : data_rom <= {16'd9908, 16'd31234};
                15'd3205 : data_rom <= {16'd9911, 16'd31233};
                15'd3206 : data_rom <= {16'd9914, 16'd31232};
                15'd3207 : data_rom <= {16'd9917, 16'd31231};
                15'd3208 : data_rom <= {16'd9920, 16'd31230};
                15'd3209 : data_rom <= {16'd9923, 16'd31229};
                15'd3210 : data_rom <= {16'd9926, 16'd31228};
                15'd3211 : data_rom <= {16'd9929, 16'd31227};
                15'd3212 : data_rom <= {16'd9932, 16'd31226};
                15'd3213 : data_rom <= {16'd9935, 16'd31225};
                15'd3214 : data_rom <= {16'd9938, 16'd31224};
                15'd3215 : data_rom <= {16'd9941, 16'd31223};
                15'd3216 : data_rom <= {16'd9944, 16'd31222};
                15'd3217 : data_rom <= {16'd9947, 16'd31221};
                15'd3218 : data_rom <= {16'd9950, 16'd31220};
                15'd3219 : data_rom <= {16'd9953, 16'd31219};
                15'd3220 : data_rom <= {16'd9956, 16'd31218};
                15'd3221 : data_rom <= {16'd9958, 16'd31217};
                15'd3222 : data_rom <= {16'd9961, 16'd31216};
                15'd3223 : data_rom <= {16'd9964, 16'd31216};
                15'd3224 : data_rom <= {16'd9967, 16'd31215};
                15'd3225 : data_rom <= {16'd9970, 16'd31214};
                15'd3226 : data_rom <= {16'd9973, 16'd31213};
                15'd3227 : data_rom <= {16'd9976, 16'd31212};
                15'd3228 : data_rom <= {16'd9979, 16'd31211};
                15'd3229 : data_rom <= {16'd9982, 16'd31210};
                15'd3230 : data_rom <= {16'd9985, 16'd31209};
                15'd3231 : data_rom <= {16'd9988, 16'd31208};
                15'd3232 : data_rom <= {16'd9991, 16'd31207};
                15'd3233 : data_rom <= {16'd9994, 16'd31206};
                15'd3234 : data_rom <= {16'd9997, 16'd31205};
                15'd3235 : data_rom <= {16'd10000, 16'd31204};
                15'd3236 : data_rom <= {16'd10003, 16'd31203};
                15'd3237 : data_rom <= {16'd10006, 16'd31202};
                15'd3238 : data_rom <= {16'd10009, 16'd31201};
                15'd3239 : data_rom <= {16'd10012, 16'd31200};
                15'd3240 : data_rom <= {16'd10015, 16'd31199};
                15'd3241 : data_rom <= {16'd10018, 16'd31198};
                15'd3242 : data_rom <= {16'd10021, 16'd31197};
                15'd3243 : data_rom <= {16'd10024, 16'd31196};
                15'd3244 : data_rom <= {16'd10027, 16'd31195};
                15'd3245 : data_rom <= {16'd10030, 16'd31194};
                15'd3246 : data_rom <= {16'd10033, 16'd31193};
                15'd3247 : data_rom <= {16'd10036, 16'd31193};
                15'd3248 : data_rom <= {16'd10039, 16'd31192};
                15'd3249 : data_rom <= {16'd10042, 16'd31191};
                15'd3250 : data_rom <= {16'd10045, 16'd31190};
                15'd3251 : data_rom <= {16'd10048, 16'd31189};
                15'd3252 : data_rom <= {16'd10051, 16'd31188};
                15'd3253 : data_rom <= {16'd10054, 16'd31187};
                15'd3254 : data_rom <= {16'd10057, 16'd31186};
                15'd3255 : data_rom <= {16'd10060, 16'd31185};
                15'd3256 : data_rom <= {16'd10063, 16'd31184};
                15'd3257 : data_rom <= {16'd10066, 16'd31183};
                15'd3258 : data_rom <= {16'd10069, 16'd31182};
                15'd3259 : data_rom <= {16'd10072, 16'd31181};
                15'd3260 : data_rom <= {16'd10075, 16'd31180};
                15'd3261 : data_rom <= {16'd10078, 16'd31179};
                15'd3262 : data_rom <= {16'd10081, 16'd31178};
                15'd3263 : data_rom <= {16'd10084, 16'd31177};
                15'd3264 : data_rom <= {16'd10087, 16'd31176};
                15'd3265 : data_rom <= {16'd10090, 16'd31175};
                15'd3266 : data_rom <= {16'd10093, 16'd31174};
                15'd3267 : data_rom <= {16'd10096, 16'd31173};
                15'd3268 : data_rom <= {16'd10099, 16'd31172};
                15'd3269 : data_rom <= {16'd10102, 16'd31171};
                15'd3270 : data_rom <= {16'd10105, 16'd31170};
                15'd3271 : data_rom <= {16'd10108, 16'd31169};
                15'd3272 : data_rom <= {16'd10111, 16'd31168};
                15'd3273 : data_rom <= {16'd10114, 16'd31167};
                15'd3274 : data_rom <= {16'd10117, 16'd31166};
                15'd3275 : data_rom <= {16'd10120, 16'd31165};
                15'd3276 : data_rom <= {16'd10123, 16'd31164};
                15'd3277 : data_rom <= {16'd10126, 16'd31164};
                15'd3278 : data_rom <= {16'd10129, 16'd31163};
                15'd3279 : data_rom <= {16'd10132, 16'd31162};
                15'd3280 : data_rom <= {16'd10135, 16'd31161};
                15'd3281 : data_rom <= {16'd10138, 16'd31160};
                15'd3282 : data_rom <= {16'd10141, 16'd31159};
                15'd3283 : data_rom <= {16'd10144, 16'd31158};
                15'd3284 : data_rom <= {16'd10147, 16'd31157};
                15'd3285 : data_rom <= {16'd10150, 16'd31156};
                15'd3286 : data_rom <= {16'd10153, 16'd31155};
                15'd3287 : data_rom <= {16'd10156, 16'd31154};
                15'd3288 : data_rom <= {16'd10159, 16'd31153};
                15'd3289 : data_rom <= {16'd10162, 16'd31152};
                15'd3290 : data_rom <= {16'd10165, 16'd31151};
                15'd3291 : data_rom <= {16'd10168, 16'd31150};
                15'd3292 : data_rom <= {16'd10171, 16'd31149};
                15'd3293 : data_rom <= {16'd10174, 16'd31148};
                15'd3294 : data_rom <= {16'd10177, 16'd31147};
                15'd3295 : data_rom <= {16'd10180, 16'd31146};
                15'd3296 : data_rom <= {16'd10183, 16'd31145};
                15'd3297 : data_rom <= {16'd10186, 16'd31144};
                15'd3298 : data_rom <= {16'd10189, 16'd31143};
                15'd3299 : data_rom <= {16'd10192, 16'd31142};
                15'd3300 : data_rom <= {16'd10195, 16'd31141};
                15'd3301 : data_rom <= {16'd10198, 16'd31140};
                15'd3302 : data_rom <= {16'd10201, 16'd31139};
                15'd3303 : data_rom <= {16'd10204, 16'd31138};
                15'd3304 : data_rom <= {16'd10207, 16'd31137};
                15'd3305 : data_rom <= {16'd10210, 16'd31136};
                15'd3306 : data_rom <= {16'd10213, 16'd31135};
                15'd3307 : data_rom <= {16'd10216, 16'd31134};
                15'd3308 : data_rom <= {16'd10219, 16'd31133};
                15'd3309 : data_rom <= {16'd10222, 16'd31132};
                15'd3310 : data_rom <= {16'd10225, 16'd31131};
                15'd3311 : data_rom <= {16'd10227, 16'd31130};
                15'd3312 : data_rom <= {16'd10230, 16'd31129};
                15'd3313 : data_rom <= {16'd10233, 16'd31128};
                15'd3314 : data_rom <= {16'd10236, 16'd31127};
                15'd3315 : data_rom <= {16'd10239, 16'd31126};
                15'd3316 : data_rom <= {16'd10242, 16'd31125};
                15'd3317 : data_rom <= {16'd10245, 16'd31124};
                15'd3318 : data_rom <= {16'd10248, 16'd31123};
                15'd3319 : data_rom <= {16'd10251, 16'd31123};
                15'd3320 : data_rom <= {16'd10254, 16'd31122};
                15'd3321 : data_rom <= {16'd10257, 16'd31121};
                15'd3322 : data_rom <= {16'd10260, 16'd31120};
                15'd3323 : data_rom <= {16'd10263, 16'd31119};
                15'd3324 : data_rom <= {16'd10266, 16'd31118};
                15'd3325 : data_rom <= {16'd10269, 16'd31117};
                15'd3326 : data_rom <= {16'd10272, 16'd31116};
                15'd3327 : data_rom <= {16'd10275, 16'd31115};
                15'd3328 : data_rom <= {16'd10278, 16'd31114};
                15'd3329 : data_rom <= {16'd10281, 16'd31113};
                15'd3330 : data_rom <= {16'd10284, 16'd31112};
                15'd3331 : data_rom <= {16'd10287, 16'd31111};
                15'd3332 : data_rom <= {16'd10290, 16'd31110};
                15'd3333 : data_rom <= {16'd10293, 16'd31109};
                15'd3334 : data_rom <= {16'd10296, 16'd31108};
                15'd3335 : data_rom <= {16'd10299, 16'd31107};
                15'd3336 : data_rom <= {16'd10302, 16'd31106};
                15'd3337 : data_rom <= {16'd10305, 16'd31105};
                15'd3338 : data_rom <= {16'd10308, 16'd31104};
                15'd3339 : data_rom <= {16'd10311, 16'd31103};
                15'd3340 : data_rom <= {16'd10314, 16'd31102};
                15'd3341 : data_rom <= {16'd10317, 16'd31101};
                15'd3342 : data_rom <= {16'd10320, 16'd31100};
                15'd3343 : data_rom <= {16'd10323, 16'd31099};
                15'd3344 : data_rom <= {16'd10326, 16'd31098};
                15'd3345 : data_rom <= {16'd10329, 16'd31097};
                15'd3346 : data_rom <= {16'd10332, 16'd31096};
                15'd3347 : data_rom <= {16'd10335, 16'd31095};
                15'd3348 : data_rom <= {16'd10338, 16'd31094};
                15'd3349 : data_rom <= {16'd10341, 16'd31093};
                15'd3350 : data_rom <= {16'd10344, 16'd31092};
                15'd3351 : data_rom <= {16'd10347, 16'd31091};
                15'd3352 : data_rom <= {16'd10350, 16'd31090};
                15'd3353 : data_rom <= {16'd10353, 16'd31089};
                15'd3354 : data_rom <= {16'd10356, 16'd31088};
                15'd3355 : data_rom <= {16'd10359, 16'd31087};
                15'd3356 : data_rom <= {16'd10362, 16'd31086};
                15'd3357 : data_rom <= {16'd10365, 16'd31085};
                15'd3358 : data_rom <= {16'd10368, 16'd31084};
                15'd3359 : data_rom <= {16'd10371, 16'd31083};
                15'd3360 : data_rom <= {16'd10374, 16'd31082};
                15'd3361 : data_rom <= {16'd10377, 16'd31081};
                15'd3362 : data_rom <= {16'd10380, 16'd31080};
                15'd3363 : data_rom <= {16'd10383, 16'd31079};
                15'd3364 : data_rom <= {16'd10386, 16'd31078};
                15'd3365 : data_rom <= {16'd10389, 16'd31077};
                15'd3366 : data_rom <= {16'd10392, 16'd31076};
                15'd3367 : data_rom <= {16'd10394, 16'd31075};
                15'd3368 : data_rom <= {16'd10397, 16'd31074};
                15'd3369 : data_rom <= {16'd10400, 16'd31073};
                15'd3370 : data_rom <= {16'd10403, 16'd31072};
                15'd3371 : data_rom <= {16'd10406, 16'd31071};
                15'd3372 : data_rom <= {16'd10409, 16'd31070};
                15'd3373 : data_rom <= {16'd10412, 16'd31069};
                15'd3374 : data_rom <= {16'd10415, 16'd31068};
                15'd3375 : data_rom <= {16'd10418, 16'd31067};
                15'd3376 : data_rom <= {16'd10421, 16'd31066};
                15'd3377 : data_rom <= {16'd10424, 16'd31065};
                15'd3378 : data_rom <= {16'd10427, 16'd31064};
                15'd3379 : data_rom <= {16'd10430, 16'd31063};
                15'd3380 : data_rom <= {16'd10433, 16'd31062};
                15'd3381 : data_rom <= {16'd10436, 16'd31061};
                15'd3382 : data_rom <= {16'd10439, 16'd31060};
                15'd3383 : data_rom <= {16'd10442, 16'd31059};
                15'd3384 : data_rom <= {16'd10445, 16'd31058};
                15'd3385 : data_rom <= {16'd10448, 16'd31057};
                15'd3386 : data_rom <= {16'd10451, 16'd31056};
                15'd3387 : data_rom <= {16'd10454, 16'd31055};
                15'd3388 : data_rom <= {16'd10457, 16'd31054};
                15'd3389 : data_rom <= {16'd10460, 16'd31053};
                15'd3390 : data_rom <= {16'd10463, 16'd31052};
                15'd3391 : data_rom <= {16'd10466, 16'd31051};
                15'd3392 : data_rom <= {16'd10469, 16'd31050};
                15'd3393 : data_rom <= {16'd10472, 16'd31049};
                15'd3394 : data_rom <= {16'd10475, 16'd31048};
                15'd3395 : data_rom <= {16'd10478, 16'd31047};
                15'd3396 : data_rom <= {16'd10481, 16'd31046};
                15'd3397 : data_rom <= {16'd10484, 16'd31045};
                15'd3398 : data_rom <= {16'd10487, 16'd31044};
                15'd3399 : data_rom <= {16'd10490, 16'd31043};
                15'd3400 : data_rom <= {16'd10493, 16'd31042};
                15'd3401 : data_rom <= {16'd10496, 16'd31041};
                15'd3402 : data_rom <= {16'd10499, 16'd31040};
                15'd3403 : data_rom <= {16'd10502, 16'd31039};
                15'd3404 : data_rom <= {16'd10505, 16'd31038};
                15'd3405 : data_rom <= {16'd10508, 16'd31037};
                15'd3406 : data_rom <= {16'd10511, 16'd31036};
                15'd3407 : data_rom <= {16'd10514, 16'd31035};
                15'd3408 : data_rom <= {16'd10517, 16'd31034};
                15'd3409 : data_rom <= {16'd10520, 16'd31033};
                15'd3410 : data_rom <= {16'd10523, 16'd31032};
                15'd3411 : data_rom <= {16'd10525, 16'd31031};
                15'd3412 : data_rom <= {16'd10528, 16'd31030};
                15'd3413 : data_rom <= {16'd10531, 16'd31029};
                15'd3414 : data_rom <= {16'd10534, 16'd31028};
                15'd3415 : data_rom <= {16'd10537, 16'd31027};
                15'd3416 : data_rom <= {16'd10540, 16'd31026};
                15'd3417 : data_rom <= {16'd10543, 16'd31025};
                15'd3418 : data_rom <= {16'd10546, 16'd31024};
                15'd3419 : data_rom <= {16'd10549, 16'd31023};
                15'd3420 : data_rom <= {16'd10552, 16'd31022};
                15'd3421 : data_rom <= {16'd10555, 16'd31021};
                15'd3422 : data_rom <= {16'd10558, 16'd31020};
                15'd3423 : data_rom <= {16'd10561, 16'd31019};
                15'd3424 : data_rom <= {16'd10564, 16'd31018};
                15'd3425 : data_rom <= {16'd10567, 16'd31017};
                15'd3426 : data_rom <= {16'd10570, 16'd31016};
                15'd3427 : data_rom <= {16'd10573, 16'd31015};
                15'd3428 : data_rom <= {16'd10576, 16'd31014};
                15'd3429 : data_rom <= {16'd10579, 16'd31013};
                15'd3430 : data_rom <= {16'd10582, 16'd31012};
                15'd3431 : data_rom <= {16'd10585, 16'd31011};
                15'd3432 : data_rom <= {16'd10588, 16'd31010};
                15'd3433 : data_rom <= {16'd10591, 16'd31009};
                15'd3434 : data_rom <= {16'd10594, 16'd31008};
                15'd3435 : data_rom <= {16'd10597, 16'd31007};
                15'd3436 : data_rom <= {16'd10600, 16'd31006};
                15'd3437 : data_rom <= {16'd10603, 16'd31005};
                15'd3438 : data_rom <= {16'd10606, 16'd31004};
                15'd3439 : data_rom <= {16'd10609, 16'd31002};
                15'd3440 : data_rom <= {16'd10612, 16'd31001};
                15'd3441 : data_rom <= {16'd10615, 16'd31000};
                15'd3442 : data_rom <= {16'd10618, 16'd30999};
                15'd3443 : data_rom <= {16'd10621, 16'd30998};
                15'd3444 : data_rom <= {16'd10624, 16'd30997};
                15'd3445 : data_rom <= {16'd10627, 16'd30996};
                15'd3446 : data_rom <= {16'd10630, 16'd30995};
                15'd3447 : data_rom <= {16'd10633, 16'd30994};
                15'd3448 : data_rom <= {16'd10635, 16'd30993};
                15'd3449 : data_rom <= {16'd10638, 16'd30992};
                15'd3450 : data_rom <= {16'd10641, 16'd30991};
                15'd3451 : data_rom <= {16'd10644, 16'd30990};
                15'd3452 : data_rom <= {16'd10647, 16'd30989};
                15'd3453 : data_rom <= {16'd10650, 16'd30988};
                15'd3454 : data_rom <= {16'd10653, 16'd30987};
                15'd3455 : data_rom <= {16'd10656, 16'd30986};
                15'd3456 : data_rom <= {16'd10659, 16'd30985};
                15'd3457 : data_rom <= {16'd10662, 16'd30984};
                15'd3458 : data_rom <= {16'd10665, 16'd30983};
                15'd3459 : data_rom <= {16'd10668, 16'd30982};
                15'd3460 : data_rom <= {16'd10671, 16'd30981};
                15'd3461 : data_rom <= {16'd10674, 16'd30980};
                15'd3462 : data_rom <= {16'd10677, 16'd30979};
                15'd3463 : data_rom <= {16'd10680, 16'd30978};
                15'd3464 : data_rom <= {16'd10683, 16'd30977};
                15'd3465 : data_rom <= {16'd10686, 16'd30976};
                15'd3466 : data_rom <= {16'd10689, 16'd30975};
                15'd3467 : data_rom <= {16'd10692, 16'd30974};
                15'd3468 : data_rom <= {16'd10695, 16'd30973};
                15'd3469 : data_rom <= {16'd10698, 16'd30972};
                15'd3470 : data_rom <= {16'd10701, 16'd30971};
                15'd3471 : data_rom <= {16'd10704, 16'd30970};
                15'd3472 : data_rom <= {16'd10707, 16'd30969};
                15'd3473 : data_rom <= {16'd10710, 16'd30968};
                15'd3474 : data_rom <= {16'd10713, 16'd30967};
                15'd3475 : data_rom <= {16'd10716, 16'd30966};
                15'd3476 : data_rom <= {16'd10719, 16'd30965};
                15'd3477 : data_rom <= {16'd10722, 16'd30964};
                15'd3478 : data_rom <= {16'd10725, 16'd30963};
                15'd3479 : data_rom <= {16'd10728, 16'd30962};
                15'd3480 : data_rom <= {16'd10731, 16'd30961};
                15'd3481 : data_rom <= {16'd10733, 16'd30960};
                15'd3482 : data_rom <= {16'd10736, 16'd30958};
                15'd3483 : data_rom <= {16'd10739, 16'd30957};
                15'd3484 : data_rom <= {16'd10742, 16'd30956};
                15'd3485 : data_rom <= {16'd10745, 16'd30955};
                15'd3486 : data_rom <= {16'd10748, 16'd30954};
                15'd3487 : data_rom <= {16'd10751, 16'd30953};
                15'd3488 : data_rom <= {16'd10754, 16'd30952};
                15'd3489 : data_rom <= {16'd10757, 16'd30951};
                15'd3490 : data_rom <= {16'd10760, 16'd30950};
                15'd3491 : data_rom <= {16'd10763, 16'd30949};
                15'd3492 : data_rom <= {16'd10766, 16'd30948};
                15'd3493 : data_rom <= {16'd10769, 16'd30947};
                15'd3494 : data_rom <= {16'd10772, 16'd30946};
                15'd3495 : data_rom <= {16'd10775, 16'd30945};
                15'd3496 : data_rom <= {16'd10778, 16'd30944};
                15'd3497 : data_rom <= {16'd10781, 16'd30943};
                15'd3498 : data_rom <= {16'd10784, 16'd30942};
                15'd3499 : data_rom <= {16'd10787, 16'd30941};
                15'd3500 : data_rom <= {16'd10790, 16'd30940};
                15'd3501 : data_rom <= {16'd10793, 16'd30939};
                15'd3502 : data_rom <= {16'd10796, 16'd30938};
                15'd3503 : data_rom <= {16'd10799, 16'd30937};
                15'd3504 : data_rom <= {16'd10802, 16'd30936};
                15'd3505 : data_rom <= {16'd10805, 16'd30935};
                15'd3506 : data_rom <= {16'd10808, 16'd30934};
                15'd3507 : data_rom <= {16'd10811, 16'd30933};
                15'd3508 : data_rom <= {16'd10814, 16'd30932};
                15'd3509 : data_rom <= {16'd10817, 16'd30931};
                15'd3510 : data_rom <= {16'd10820, 16'd30930};
                15'd3511 : data_rom <= {16'd10822, 16'd30929};
                15'd3512 : data_rom <= {16'd10825, 16'd30927};
                15'd3513 : data_rom <= {16'd10828, 16'd30926};
                15'd3514 : data_rom <= {16'd10831, 16'd30925};
                15'd3515 : data_rom <= {16'd10834, 16'd30924};
                15'd3516 : data_rom <= {16'd10837, 16'd30923};
                15'd3517 : data_rom <= {16'd10840, 16'd30922};
                15'd3518 : data_rom <= {16'd10843, 16'd30921};
                15'd3519 : data_rom <= {16'd10846, 16'd30920};
                15'd3520 : data_rom <= {16'd10849, 16'd30919};
                15'd3521 : data_rom <= {16'd10852, 16'd30918};
                15'd3522 : data_rom <= {16'd10855, 16'd30917};
                15'd3523 : data_rom <= {16'd10858, 16'd30916};
                15'd3524 : data_rom <= {16'd10861, 16'd30915};
                15'd3525 : data_rom <= {16'd10864, 16'd30914};
                15'd3526 : data_rom <= {16'd10867, 16'd30913};
                15'd3527 : data_rom <= {16'd10870, 16'd30912};
                15'd3528 : data_rom <= {16'd10873, 16'd30911};
                15'd3529 : data_rom <= {16'd10876, 16'd30910};
                15'd3530 : data_rom <= {16'd10879, 16'd30909};
                15'd3531 : data_rom <= {16'd10882, 16'd30908};
                15'd3532 : data_rom <= {16'd10885, 16'd30907};
                15'd3533 : data_rom <= {16'd10888, 16'd30906};
                15'd3534 : data_rom <= {16'd10891, 16'd30905};
                15'd3535 : data_rom <= {16'd10894, 16'd30904};
                15'd3536 : data_rom <= {16'd10897, 16'd30902};
                15'd3537 : data_rom <= {16'd10900, 16'd30901};
                15'd3538 : data_rom <= {16'd10903, 16'd30900};
                15'd3539 : data_rom <= {16'd10905, 16'd30899};
                15'd3540 : data_rom <= {16'd10908, 16'd30898};
                15'd3541 : data_rom <= {16'd10911, 16'd30897};
                15'd3542 : data_rom <= {16'd10914, 16'd30896};
                15'd3543 : data_rom <= {16'd10917, 16'd30895};
                15'd3544 : data_rom <= {16'd10920, 16'd30894};
                15'd3545 : data_rom <= {16'd10923, 16'd30893};
                15'd3546 : data_rom <= {16'd10926, 16'd30892};
                15'd3547 : data_rom <= {16'd10929, 16'd30891};
                15'd3548 : data_rom <= {16'd10932, 16'd30890};
                15'd3549 : data_rom <= {16'd10935, 16'd30889};
                15'd3550 : data_rom <= {16'd10938, 16'd30888};
                15'd3551 : data_rom <= {16'd10941, 16'd30887};
                15'd3552 : data_rom <= {16'd10944, 16'd30886};
                15'd3553 : data_rom <= {16'd10947, 16'd30885};
                15'd3554 : data_rom <= {16'd10950, 16'd30884};
                15'd3555 : data_rom <= {16'd10953, 16'd30883};
                15'd3556 : data_rom <= {16'd10956, 16'd30882};
                15'd3557 : data_rom <= {16'd10959, 16'd30880};
                15'd3558 : data_rom <= {16'd10962, 16'd30879};
                15'd3559 : data_rom <= {16'd10965, 16'd30878};
                15'd3560 : data_rom <= {16'd10968, 16'd30877};
                15'd3561 : data_rom <= {16'd10971, 16'd30876};
                15'd3562 : data_rom <= {16'd10974, 16'd30875};
                15'd3563 : data_rom <= {16'd10977, 16'd30874};
                15'd3564 : data_rom <= {16'd10980, 16'd30873};
                15'd3565 : data_rom <= {16'd10982, 16'd30872};
                15'd3566 : data_rom <= {16'd10985, 16'd30871};
                15'd3567 : data_rom <= {16'd10988, 16'd30870};
                15'd3568 : data_rom <= {16'd10991, 16'd30869};
                15'd3569 : data_rom <= {16'd10994, 16'd30868};
                15'd3570 : data_rom <= {16'd10997, 16'd30867};
                15'd3571 : data_rom <= {16'd11000, 16'd30866};
                15'd3572 : data_rom <= {16'd11003, 16'd30865};
                15'd3573 : data_rom <= {16'd11006, 16'd30864};
                15'd3574 : data_rom <= {16'd11009, 16'd30863};
                15'd3575 : data_rom <= {16'd11012, 16'd30862};
                15'd3576 : data_rom <= {16'd11015, 16'd30860};
                15'd3577 : data_rom <= {16'd11018, 16'd30859};
                15'd3578 : data_rom <= {16'd11021, 16'd30858};
                15'd3579 : data_rom <= {16'd11024, 16'd30857};
                15'd3580 : data_rom <= {16'd11027, 16'd30856};
                15'd3581 : data_rom <= {16'd11030, 16'd30855};
                15'd3582 : data_rom <= {16'd11033, 16'd30854};
                15'd3583 : data_rom <= {16'd11036, 16'd30853};
                15'd3584 : data_rom <= {16'd11039, 16'd30852};
                15'd3585 : data_rom <= {16'd11042, 16'd30851};
                15'd3586 : data_rom <= {16'd11045, 16'd30850};
                15'd3587 : data_rom <= {16'd11048, 16'd30849};
                15'd3588 : data_rom <= {16'd11051, 16'd30848};
                15'd3589 : data_rom <= {16'd11053, 16'd30847};
                15'd3590 : data_rom <= {16'd11056, 16'd30846};
                15'd3591 : data_rom <= {16'd11059, 16'd30845};
                15'd3592 : data_rom <= {16'd11062, 16'd30844};
                15'd3593 : data_rom <= {16'd11065, 16'd30842};
                15'd3594 : data_rom <= {16'd11068, 16'd30841};
                15'd3595 : data_rom <= {16'd11071, 16'd30840};
                15'd3596 : data_rom <= {16'd11074, 16'd30839};
                15'd3597 : data_rom <= {16'd11077, 16'd30838};
                15'd3598 : data_rom <= {16'd11080, 16'd30837};
                15'd3599 : data_rom <= {16'd11083, 16'd30836};
                15'd3600 : data_rom <= {16'd11086, 16'd30835};
                15'd3601 : data_rom <= {16'd11089, 16'd30834};
                15'd3602 : data_rom <= {16'd11092, 16'd30833};
                15'd3603 : data_rom <= {16'd11095, 16'd30832};
                15'd3604 : data_rom <= {16'd11098, 16'd30831};
                15'd3605 : data_rom <= {16'd11101, 16'd30830};
                15'd3606 : data_rom <= {16'd11104, 16'd30829};
                15'd3607 : data_rom <= {16'd11107, 16'd30828};
                15'd3608 : data_rom <= {16'd11110, 16'd30827};
                15'd3609 : data_rom <= {16'd11113, 16'd30825};
                15'd3610 : data_rom <= {16'd11116, 16'd30824};
                15'd3611 : data_rom <= {16'd11119, 16'd30823};
                15'd3612 : data_rom <= {16'd11121, 16'd30822};
                15'd3613 : data_rom <= {16'd11124, 16'd30821};
                15'd3614 : data_rom <= {16'd11127, 16'd30820};
                15'd3615 : data_rom <= {16'd11130, 16'd30819};
                15'd3616 : data_rom <= {16'd11133, 16'd30818};
                15'd3617 : data_rom <= {16'd11136, 16'd30817};
                15'd3618 : data_rom <= {16'd11139, 16'd30816};
                15'd3619 : data_rom <= {16'd11142, 16'd30815};
                15'd3620 : data_rom <= {16'd11145, 16'd30814};
                15'd3621 : data_rom <= {16'd11148, 16'd30813};
                15'd3622 : data_rom <= {16'd11151, 16'd30812};
                15'd3623 : data_rom <= {16'd11154, 16'd30811};
                15'd3624 : data_rom <= {16'd11157, 16'd30809};
                15'd3625 : data_rom <= {16'd11160, 16'd30808};
                15'd3626 : data_rom <= {16'd11163, 16'd30807};
                15'd3627 : data_rom <= {16'd11166, 16'd30806};
                15'd3628 : data_rom <= {16'd11169, 16'd30805};
                15'd3629 : data_rom <= {16'd11172, 16'd30804};
                15'd3630 : data_rom <= {16'd11175, 16'd30803};
                15'd3631 : data_rom <= {16'd11178, 16'd30802};
                15'd3632 : data_rom <= {16'd11181, 16'd30801};
                15'd3633 : data_rom <= {16'd11184, 16'd30800};
                15'd3634 : data_rom <= {16'd11186, 16'd30799};
                15'd3635 : data_rom <= {16'd11189, 16'd30798};
                15'd3636 : data_rom <= {16'd11192, 16'd30797};
                15'd3637 : data_rom <= {16'd11195, 16'd30796};
                15'd3638 : data_rom <= {16'd11198, 16'd30794};
                15'd3639 : data_rom <= {16'd11201, 16'd30793};
                15'd3640 : data_rom <= {16'd11204, 16'd30792};
                15'd3641 : data_rom <= {16'd11207, 16'd30791};
                15'd3642 : data_rom <= {16'd11210, 16'd30790};
                15'd3643 : data_rom <= {16'd11213, 16'd30789};
                15'd3644 : data_rom <= {16'd11216, 16'd30788};
                15'd3645 : data_rom <= {16'd11219, 16'd30787};
                15'd3646 : data_rom <= {16'd11222, 16'd30786};
                15'd3647 : data_rom <= {16'd11225, 16'd30785};
                15'd3648 : data_rom <= {16'd11228, 16'd30784};
                15'd3649 : data_rom <= {16'd11231, 16'd30783};
                15'd3650 : data_rom <= {16'd11234, 16'd30782};
                15'd3651 : data_rom <= {16'd11237, 16'd30780};
                15'd3652 : data_rom <= {16'd11240, 16'd30779};
                15'd3653 : data_rom <= {16'd11243, 16'd30778};
                15'd3654 : data_rom <= {16'd11246, 16'd30777};
                15'd3655 : data_rom <= {16'd11248, 16'd30776};
                15'd3656 : data_rom <= {16'd11251, 16'd30775};
                15'd3657 : data_rom <= {16'd11254, 16'd30774};
                15'd3658 : data_rom <= {16'd11257, 16'd30773};
                15'd3659 : data_rom <= {16'd11260, 16'd30772};
                15'd3660 : data_rom <= {16'd11263, 16'd30771};
                15'd3661 : data_rom <= {16'd11266, 16'd30770};
                15'd3662 : data_rom <= {16'd11269, 16'd30769};
                15'd3663 : data_rom <= {16'd11272, 16'd30768};
                15'd3664 : data_rom <= {16'd11275, 16'd30766};
                15'd3665 : data_rom <= {16'd11278, 16'd30765};
                15'd3666 : data_rom <= {16'd11281, 16'd30764};
                15'd3667 : data_rom <= {16'd11284, 16'd30763};
                15'd3668 : data_rom <= {16'd11287, 16'd30762};
                15'd3669 : data_rom <= {16'd11290, 16'd30761};
                15'd3670 : data_rom <= {16'd11293, 16'd30760};
                15'd3671 : data_rom <= {16'd11296, 16'd30759};
                15'd3672 : data_rom <= {16'd11299, 16'd30758};
                15'd3673 : data_rom <= {16'd11302, 16'd30757};
                15'd3674 : data_rom <= {16'd11304, 16'd30756};
                15'd3675 : data_rom <= {16'd11307, 16'd30755};
                15'd3676 : data_rom <= {16'd11310, 16'd30753};
                15'd3677 : data_rom <= {16'd11313, 16'd30752};
                15'd3678 : data_rom <= {16'd11316, 16'd30751};
                15'd3679 : data_rom <= {16'd11319, 16'd30750};
                15'd3680 : data_rom <= {16'd11322, 16'd30749};
                15'd3681 : data_rom <= {16'd11325, 16'd30748};
                15'd3682 : data_rom <= {16'd11328, 16'd30747};
                15'd3683 : data_rom <= {16'd11331, 16'd30746};
                15'd3684 : data_rom <= {16'd11334, 16'd30745};
                15'd3685 : data_rom <= {16'd11337, 16'd30744};
                15'd3686 : data_rom <= {16'd11340, 16'd30743};
                15'd3687 : data_rom <= {16'd11343, 16'd30742};
                15'd3688 : data_rom <= {16'd11346, 16'd30740};
                15'd3689 : data_rom <= {16'd11349, 16'd30739};
                15'd3690 : data_rom <= {16'd11352, 16'd30738};
                15'd3691 : data_rom <= {16'd11355, 16'd30737};
                15'd3692 : data_rom <= {16'd11358, 16'd30736};
                15'd3693 : data_rom <= {16'd11361, 16'd30735};
                15'd3694 : data_rom <= {16'd11363, 16'd30734};
                15'd3695 : data_rom <= {16'd11366, 16'd30733};
                15'd3696 : data_rom <= {16'd11369, 16'd30732};
                15'd3697 : data_rom <= {16'd11372, 16'd30731};
                15'd3698 : data_rom <= {16'd11375, 16'd30730};
                15'd3699 : data_rom <= {16'd11378, 16'd30728};
                15'd3700 : data_rom <= {16'd11381, 16'd30727};
                15'd3701 : data_rom <= {16'd11384, 16'd30726};
                15'd3702 : data_rom <= {16'd11387, 16'd30725};
                15'd3703 : data_rom <= {16'd11390, 16'd30724};
                15'd3704 : data_rom <= {16'd11393, 16'd30723};
                15'd3705 : data_rom <= {16'd11396, 16'd30722};
                15'd3706 : data_rom <= {16'd11399, 16'd30721};
                15'd3707 : data_rom <= {16'd11402, 16'd30720};
                15'd3708 : data_rom <= {16'd11405, 16'd30719};
                15'd3709 : data_rom <= {16'd11408, 16'd30718};
                15'd3710 : data_rom <= {16'd11411, 16'd30716};
                15'd3711 : data_rom <= {16'd11414, 16'd30715};
                15'd3712 : data_rom <= {16'd11416, 16'd30714};
                15'd3713 : data_rom <= {16'd11419, 16'd30713};
                15'd3714 : data_rom <= {16'd11422, 16'd30712};
                15'd3715 : data_rom <= {16'd11425, 16'd30711};
                15'd3716 : data_rom <= {16'd11428, 16'd30710};
                15'd3717 : data_rom <= {16'd11431, 16'd30709};
                15'd3718 : data_rom <= {16'd11434, 16'd30708};
                15'd3719 : data_rom <= {16'd11437, 16'd30707};
                15'd3720 : data_rom <= {16'd11440, 16'd30705};
                15'd3721 : data_rom <= {16'd11443, 16'd30704};
                15'd3722 : data_rom <= {16'd11446, 16'd30703};
                15'd3723 : data_rom <= {16'd11449, 16'd30702};
                15'd3724 : data_rom <= {16'd11452, 16'd30701};
                15'd3725 : data_rom <= {16'd11455, 16'd30700};
                15'd3726 : data_rom <= {16'd11458, 16'd30699};
                15'd3727 : data_rom <= {16'd11461, 16'd30698};
                15'd3728 : data_rom <= {16'd11464, 16'd30697};
                15'd3729 : data_rom <= {16'd11467, 16'd30696};
                15'd3730 : data_rom <= {16'd11469, 16'd30694};
                15'd3731 : data_rom <= {16'd11472, 16'd30693};
                15'd3732 : data_rom <= {16'd11475, 16'd30692};
                15'd3733 : data_rom <= {16'd11478, 16'd30691};
                15'd3734 : data_rom <= {16'd11481, 16'd30690};
                15'd3735 : data_rom <= {16'd11484, 16'd30689};
                15'd3736 : data_rom <= {16'd11487, 16'd30688};
                15'd3737 : data_rom <= {16'd11490, 16'd30687};
                15'd3738 : data_rom <= {16'd11493, 16'd30686};
                15'd3739 : data_rom <= {16'd11496, 16'd30685};
                15'd3740 : data_rom <= {16'd11499, 16'd30683};
                15'd3741 : data_rom <= {16'd11502, 16'd30682};
                15'd3742 : data_rom <= {16'd11505, 16'd30681};
                15'd3743 : data_rom <= {16'd11508, 16'd30680};
                15'd3744 : data_rom <= {16'd11511, 16'd30679};
                15'd3745 : data_rom <= {16'd11514, 16'd30678};
                15'd3746 : data_rom <= {16'd11517, 16'd30677};
                15'd3747 : data_rom <= {16'd11519, 16'd30676};
                15'd3748 : data_rom <= {16'd11522, 16'd30675};
                15'd3749 : data_rom <= {16'd11525, 16'd30674};
                15'd3750 : data_rom <= {16'd11528, 16'd30672};
                15'd3751 : data_rom <= {16'd11531, 16'd30671};
                15'd3752 : data_rom <= {16'd11534, 16'd30670};
                15'd3753 : data_rom <= {16'd11537, 16'd30669};
                15'd3754 : data_rom <= {16'd11540, 16'd30668};
                15'd3755 : data_rom <= {16'd11543, 16'd30667};
                15'd3756 : data_rom <= {16'd11546, 16'd30666};
                15'd3757 : data_rom <= {16'd11549, 16'd30665};
                15'd3758 : data_rom <= {16'd11552, 16'd30664};
                15'd3759 : data_rom <= {16'd11555, 16'd30662};
                15'd3760 : data_rom <= {16'd11558, 16'd30661};
                15'd3761 : data_rom <= {16'd11561, 16'd30660};
                15'd3762 : data_rom <= {16'd11564, 16'd30659};
                15'd3763 : data_rom <= {16'd11567, 16'd30658};
                15'd3764 : data_rom <= {16'd11569, 16'd30657};
                15'd3765 : data_rom <= {16'd11572, 16'd30656};
                15'd3766 : data_rom <= {16'd11575, 16'd30655};
                15'd3767 : data_rom <= {16'd11578, 16'd30654};
                15'd3768 : data_rom <= {16'd11581, 16'd30652};
                15'd3769 : data_rom <= {16'd11584, 16'd30651};
                15'd3770 : data_rom <= {16'd11587, 16'd30650};
                15'd3771 : data_rom <= {16'd11590, 16'd30649};
                15'd3772 : data_rom <= {16'd11593, 16'd30648};
                15'd3773 : data_rom <= {16'd11596, 16'd30647};
                15'd3774 : data_rom <= {16'd11599, 16'd30646};
                15'd3775 : data_rom <= {16'd11602, 16'd30645};
                15'd3776 : data_rom <= {16'd11605, 16'd30644};
                15'd3777 : data_rom <= {16'd11608, 16'd30642};
                15'd3778 : data_rom <= {16'd11611, 16'd30641};
                15'd3779 : data_rom <= {16'd11614, 16'd30640};
                15'd3780 : data_rom <= {16'd11616, 16'd30639};
                15'd3781 : data_rom <= {16'd11619, 16'd30638};
                15'd3782 : data_rom <= {16'd11622, 16'd30637};
                15'd3783 : data_rom <= {16'd11625, 16'd30636};
                15'd3784 : data_rom <= {16'd11628, 16'd30635};
                15'd3785 : data_rom <= {16'd11631, 16'd30634};
                15'd3786 : data_rom <= {16'd11634, 16'd30632};
                15'd3787 : data_rom <= {16'd11637, 16'd30631};
                15'd3788 : data_rom <= {16'd11640, 16'd30630};
                15'd3789 : data_rom <= {16'd11643, 16'd30629};
                15'd3790 : data_rom <= {16'd11646, 16'd30628};
                15'd3791 : data_rom <= {16'd11649, 16'd30627};
                15'd3792 : data_rom <= {16'd11652, 16'd30626};
                15'd3793 : data_rom <= {16'd11655, 16'd30625};
                15'd3794 : data_rom <= {16'd11658, 16'd30624};
                15'd3795 : data_rom <= {16'd11661, 16'd30622};
                15'd3796 : data_rom <= {16'd11663, 16'd30621};
                15'd3797 : data_rom <= {16'd11666, 16'd30620};
                15'd3798 : data_rom <= {16'd11669, 16'd30619};
                15'd3799 : data_rom <= {16'd11672, 16'd30618};
                15'd3800 : data_rom <= {16'd11675, 16'd30617};
                15'd3801 : data_rom <= {16'd11678, 16'd30616};
                15'd3802 : data_rom <= {16'd11681, 16'd30615};
                15'd3803 : data_rom <= {16'd11684, 16'd30613};
                15'd3804 : data_rom <= {16'd11687, 16'd30612};
                15'd3805 : data_rom <= {16'd11690, 16'd30611};
                15'd3806 : data_rom <= {16'd11693, 16'd30610};
                15'd3807 : data_rom <= {16'd11696, 16'd30609};
                15'd3808 : data_rom <= {16'd11699, 16'd30608};
                15'd3809 : data_rom <= {16'd11702, 16'd30607};
                15'd3810 : data_rom <= {16'd11705, 16'd30606};
                15'd3811 : data_rom <= {16'd11707, 16'd30604};
                15'd3812 : data_rom <= {16'd11710, 16'd30603};
                15'd3813 : data_rom <= {16'd11713, 16'd30602};
                15'd3814 : data_rom <= {16'd11716, 16'd30601};
                15'd3815 : data_rom <= {16'd11719, 16'd30600};
                15'd3816 : data_rom <= {16'd11722, 16'd30599};
                15'd3817 : data_rom <= {16'd11725, 16'd30598};
                15'd3818 : data_rom <= {16'd11728, 16'd30597};
                15'd3819 : data_rom <= {16'd11731, 16'd30595};
                15'd3820 : data_rom <= {16'd11734, 16'd30594};
                15'd3821 : data_rom <= {16'd11737, 16'd30593};
                15'd3822 : data_rom <= {16'd11740, 16'd30592};
                15'd3823 : data_rom <= {16'd11743, 16'd30591};
                15'd3824 : data_rom <= {16'd11746, 16'd30590};
                15'd3825 : data_rom <= {16'd11749, 16'd30589};
                15'd3826 : data_rom <= {16'd11751, 16'd30588};
                15'd3827 : data_rom <= {16'd11754, 16'd30586};
                15'd3828 : data_rom <= {16'd11757, 16'd30585};
                15'd3829 : data_rom <= {16'd11760, 16'd30584};
                15'd3830 : data_rom <= {16'd11763, 16'd30583};
                15'd3831 : data_rom <= {16'd11766, 16'd30582};
                15'd3832 : data_rom <= {16'd11769, 16'd30581};
                15'd3833 : data_rom <= {16'd11772, 16'd30580};
                15'd3834 : data_rom <= {16'd11775, 16'd30579};
                15'd3835 : data_rom <= {16'd11778, 16'd30577};
                15'd3836 : data_rom <= {16'd11781, 16'd30576};
                15'd3837 : data_rom <= {16'd11784, 16'd30575};
                15'd3838 : data_rom <= {16'd11787, 16'd30574};
                15'd3839 : data_rom <= {16'd11790, 16'd30573};
                15'd3840 : data_rom <= {16'd11793, 16'd30572};
                15'd3841 : data_rom <= {16'd11795, 16'd30571};
                15'd3842 : data_rom <= {16'd11798, 16'd30570};
                15'd3843 : data_rom <= {16'd11801, 16'd30568};
                15'd3844 : data_rom <= {16'd11804, 16'd30567};
                15'd3845 : data_rom <= {16'd11807, 16'd30566};
                15'd3846 : data_rom <= {16'd11810, 16'd30565};
                15'd3847 : data_rom <= {16'd11813, 16'd30564};
                15'd3848 : data_rom <= {16'd11816, 16'd30563};
                15'd3849 : data_rom <= {16'd11819, 16'd30562};
                15'd3850 : data_rom <= {16'd11822, 16'd30560};
                15'd3851 : data_rom <= {16'd11825, 16'd30559};
                15'd3852 : data_rom <= {16'd11828, 16'd30558};
                15'd3853 : data_rom <= {16'd11831, 16'd30557};
                15'd3854 : data_rom <= {16'd11834, 16'd30556};
                15'd3855 : data_rom <= {16'd11836, 16'd30555};
                15'd3856 : data_rom <= {16'd11839, 16'd30554};
                15'd3857 : data_rom <= {16'd11842, 16'd30553};
                15'd3858 : data_rom <= {16'd11845, 16'd30551};
                15'd3859 : data_rom <= {16'd11848, 16'd30550};
                15'd3860 : data_rom <= {16'd11851, 16'd30549};
                15'd3861 : data_rom <= {16'd11854, 16'd30548};
                15'd3862 : data_rom <= {16'd11857, 16'd30547};
                15'd3863 : data_rom <= {16'd11860, 16'd30546};
                15'd3864 : data_rom <= {16'd11863, 16'd30545};
                15'd3865 : data_rom <= {16'd11866, 16'd30543};
                15'd3866 : data_rom <= {16'd11869, 16'd30542};
                15'd3867 : data_rom <= {16'd11872, 16'd30541};
                15'd3868 : data_rom <= {16'd11875, 16'd30540};
                15'd3869 : data_rom <= {16'd11877, 16'd30539};
                15'd3870 : data_rom <= {16'd11880, 16'd30538};
                15'd3871 : data_rom <= {16'd11883, 16'd30537};
                15'd3872 : data_rom <= {16'd11886, 16'd30535};
                15'd3873 : data_rom <= {16'd11889, 16'd30534};
                15'd3874 : data_rom <= {16'd11892, 16'd30533};
                15'd3875 : data_rom <= {16'd11895, 16'd30532};
                15'd3876 : data_rom <= {16'd11898, 16'd30531};
                15'd3877 : data_rom <= {16'd11901, 16'd30530};
                15'd3878 : data_rom <= {16'd11904, 16'd30529};
                15'd3879 : data_rom <= {16'd11907, 16'd30528};
                15'd3880 : data_rom <= {16'd11910, 16'd30526};
                15'd3881 : data_rom <= {16'd11913, 16'd30525};
                15'd3882 : data_rom <= {16'd11916, 16'd30524};
                15'd3883 : data_rom <= {16'd11918, 16'd30523};
                15'd3884 : data_rom <= {16'd11921, 16'd30522};
                15'd3885 : data_rom <= {16'd11924, 16'd30521};
                15'd3886 : data_rom <= {16'd11927, 16'd30520};
                15'd3887 : data_rom <= {16'd11930, 16'd30518};
                15'd3888 : data_rom <= {16'd11933, 16'd30517};
                15'd3889 : data_rom <= {16'd11936, 16'd30516};
                15'd3890 : data_rom <= {16'd11939, 16'd30515};
                15'd3891 : data_rom <= {16'd11942, 16'd30514};
                15'd3892 : data_rom <= {16'd11945, 16'd30513};
                15'd3893 : data_rom <= {16'd11948, 16'd30511};
                15'd3894 : data_rom <= {16'd11951, 16'd30510};
                15'd3895 : data_rom <= {16'd11954, 16'd30509};
                15'd3896 : data_rom <= {16'd11956, 16'd30508};
                15'd3897 : data_rom <= {16'd11959, 16'd30507};
                15'd3898 : data_rom <= {16'd11962, 16'd30506};
                15'd3899 : data_rom <= {16'd11965, 16'd30505};
                15'd3900 : data_rom <= {16'd11968, 16'd30503};
                15'd3901 : data_rom <= {16'd11971, 16'd30502};
                15'd3902 : data_rom <= {16'd11974, 16'd30501};
                15'd3903 : data_rom <= {16'd11977, 16'd30500};
                15'd3904 : data_rom <= {16'd11980, 16'd30499};
                15'd3905 : data_rom <= {16'd11983, 16'd30498};
                15'd3906 : data_rom <= {16'd11986, 16'd30497};
                15'd3907 : data_rom <= {16'd11989, 16'd30495};
                15'd3908 : data_rom <= {16'd11992, 16'd30494};
                15'd3909 : data_rom <= {16'd11995, 16'd30493};
                15'd3910 : data_rom <= {16'd11997, 16'd30492};
                15'd3911 : data_rom <= {16'd12000, 16'd30491};
                15'd3912 : data_rom <= {16'd12003, 16'd30490};
                15'd3913 : data_rom <= {16'd12006, 16'd30489};
                15'd3914 : data_rom <= {16'd12009, 16'd30487};
                15'd3915 : data_rom <= {16'd12012, 16'd30486};
                15'd3916 : data_rom <= {16'd12015, 16'd30485};
                15'd3917 : data_rom <= {16'd12018, 16'd30484};
                15'd3918 : data_rom <= {16'd12021, 16'd30483};
                15'd3919 : data_rom <= {16'd12024, 16'd30482};
                15'd3920 : data_rom <= {16'd12027, 16'd30480};
                15'd3921 : data_rom <= {16'd12030, 16'd30479};
                15'd3922 : data_rom <= {16'd12033, 16'd30478};
                15'd3923 : data_rom <= {16'd12035, 16'd30477};
                15'd3924 : data_rom <= {16'd12038, 16'd30476};
                15'd3925 : data_rom <= {16'd12041, 16'd30475};
                15'd3926 : data_rom <= {16'd12044, 16'd30474};
                15'd3927 : data_rom <= {16'd12047, 16'd30472};
                15'd3928 : data_rom <= {16'd12050, 16'd30471};
                15'd3929 : data_rom <= {16'd12053, 16'd30470};
                15'd3930 : data_rom <= {16'd12056, 16'd30469};
                15'd3931 : data_rom <= {16'd12059, 16'd30468};
                15'd3932 : data_rom <= {16'd12062, 16'd30467};
                15'd3933 : data_rom <= {16'd12065, 16'd30465};
                15'd3934 : data_rom <= {16'd12068, 16'd30464};
                15'd3935 : data_rom <= {16'd12070, 16'd30463};
                15'd3936 : data_rom <= {16'd12073, 16'd30462};
                15'd3937 : data_rom <= {16'd12076, 16'd30461};
                15'd3938 : data_rom <= {16'd12079, 16'd30460};
                15'd3939 : data_rom <= {16'd12082, 16'd30459};
                15'd3940 : data_rom <= {16'd12085, 16'd30457};
                15'd3941 : data_rom <= {16'd12088, 16'd30456};
                15'd3942 : data_rom <= {16'd12091, 16'd30455};
                15'd3943 : data_rom <= {16'd12094, 16'd30454};
                15'd3944 : data_rom <= {16'd12097, 16'd30453};
                15'd3945 : data_rom <= {16'd12100, 16'd30452};
                15'd3946 : data_rom <= {16'd12103, 16'd30450};
                15'd3947 : data_rom <= {16'd12106, 16'd30449};
                15'd3948 : data_rom <= {16'd12108, 16'd30448};
                15'd3949 : data_rom <= {16'd12111, 16'd30447};
                15'd3950 : data_rom <= {16'd12114, 16'd30446};
                15'd3951 : data_rom <= {16'd12117, 16'd30445};
                15'd3952 : data_rom <= {16'd12120, 16'd30443};
                15'd3953 : data_rom <= {16'd12123, 16'd30442};
                15'd3954 : data_rom <= {16'd12126, 16'd30441};
                15'd3955 : data_rom <= {16'd12129, 16'd30440};
                15'd3956 : data_rom <= {16'd12132, 16'd30439};
                15'd3957 : data_rom <= {16'd12135, 16'd30438};
                15'd3958 : data_rom <= {16'd12138, 16'd30436};
                15'd3959 : data_rom <= {16'd12141, 16'd30435};
                15'd3960 : data_rom <= {16'd12143, 16'd30434};
                15'd3961 : data_rom <= {16'd12146, 16'd30433};
                15'd3962 : data_rom <= {16'd12149, 16'd30432};
                15'd3963 : data_rom <= {16'd12152, 16'd30431};
                15'd3964 : data_rom <= {16'd12155, 16'd30429};
                15'd3965 : data_rom <= {16'd12158, 16'd30428};
                15'd3966 : data_rom <= {16'd12161, 16'd30427};
                15'd3967 : data_rom <= {16'd12164, 16'd30426};
                15'd3968 : data_rom <= {16'd12167, 16'd30425};
                15'd3969 : data_rom <= {16'd12170, 16'd30424};
                15'd3970 : data_rom <= {16'd12173, 16'd30422};
                15'd3971 : data_rom <= {16'd12176, 16'd30421};
                15'd3972 : data_rom <= {16'd12178, 16'd30420};
                15'd3973 : data_rom <= {16'd12181, 16'd30419};
                15'd3974 : data_rom <= {16'd12184, 16'd30418};
                15'd3975 : data_rom <= {16'd12187, 16'd30417};
                15'd3976 : data_rom <= {16'd12190, 16'd30415};
                15'd3977 : data_rom <= {16'd12193, 16'd30414};
                15'd3978 : data_rom <= {16'd12196, 16'd30413};
                15'd3979 : data_rom <= {16'd12199, 16'd30412};
                15'd3980 : data_rom <= {16'd12202, 16'd30411};
                15'd3981 : data_rom <= {16'd12205, 16'd30410};
                15'd3982 : data_rom <= {16'd12208, 16'd30408};
                15'd3983 : data_rom <= {16'd12211, 16'd30407};
                15'd3984 : data_rom <= {16'd12213, 16'd30406};
                15'd3985 : data_rom <= {16'd12216, 16'd30405};
                15'd3986 : data_rom <= {16'd12219, 16'd30404};
                15'd3987 : data_rom <= {16'd12222, 16'd30403};
                15'd3988 : data_rom <= {16'd12225, 16'd30401};
                15'd3989 : data_rom <= {16'd12228, 16'd30400};
                15'd3990 : data_rom <= {16'd12231, 16'd30399};
                15'd3991 : data_rom <= {16'd12234, 16'd30398};
                15'd3992 : data_rom <= {16'd12237, 16'd30397};
                15'd3993 : data_rom <= {16'd12240, 16'd30396};
                15'd3994 : data_rom <= {16'd12243, 16'd30394};
                15'd3995 : data_rom <= {16'd12246, 16'd30393};
                15'd3996 : data_rom <= {16'd12248, 16'd30392};
                15'd3997 : data_rom <= {16'd12251, 16'd30391};
                15'd3998 : data_rom <= {16'd12254, 16'd30390};
                15'd3999 : data_rom <= {16'd12257, 16'd30388};
                15'd4000 : data_rom <= {16'd12260, 16'd30387};
                15'd4001 : data_rom <= {16'd12263, 16'd30386};
                15'd4002 : data_rom <= {16'd12266, 16'd30385};
                15'd4003 : data_rom <= {16'd12269, 16'd30384};
                15'd4004 : data_rom <= {16'd12272, 16'd30383};
                15'd4005 : data_rom <= {16'd12275, 16'd30381};
                15'd4006 : data_rom <= {16'd12278, 16'd30380};
                15'd4007 : data_rom <= {16'd12280, 16'd30379};
                15'd4008 : data_rom <= {16'd12283, 16'd30378};
                15'd4009 : data_rom <= {16'd12286, 16'd30377};
                15'd4010 : data_rom <= {16'd12289, 16'd30376};
                15'd4011 : data_rom <= {16'd12292, 16'd30374};
                15'd4012 : data_rom <= {16'd12295, 16'd30373};
                15'd4013 : data_rom <= {16'd12298, 16'd30372};
                15'd4014 : data_rom <= {16'd12301, 16'd30371};
                15'd4015 : data_rom <= {16'd12304, 16'd30370};
                15'd4016 : data_rom <= {16'd12307, 16'd30368};
                15'd4017 : data_rom <= {16'd12310, 16'd30367};
                15'd4018 : data_rom <= {16'd12313, 16'd30366};
                15'd4019 : data_rom <= {16'd12315, 16'd30365};
                15'd4020 : data_rom <= {16'd12318, 16'd30364};
                15'd4021 : data_rom <= {16'd12321, 16'd30363};
                15'd4022 : data_rom <= {16'd12324, 16'd30361};
                15'd4023 : data_rom <= {16'd12327, 16'd30360};
                15'd4024 : data_rom <= {16'd12330, 16'd30359};
                15'd4025 : data_rom <= {16'd12333, 16'd30358};
                15'd4026 : data_rom <= {16'd12336, 16'd30357};
                15'd4027 : data_rom <= {16'd12339, 16'd30355};
                15'd4028 : data_rom <= {16'd12342, 16'd30354};
                15'd4029 : data_rom <= {16'd12345, 16'd30353};
                15'd4030 : data_rom <= {16'd12347, 16'd30352};
                15'd4031 : data_rom <= {16'd12350, 16'd30351};
                15'd4032 : data_rom <= {16'd12353, 16'd30350};
                15'd4033 : data_rom <= {16'd12356, 16'd30348};
                15'd4034 : data_rom <= {16'd12359, 16'd30347};
                15'd4035 : data_rom <= {16'd12362, 16'd30346};
                15'd4036 : data_rom <= {16'd12365, 16'd30345};
                15'd4037 : data_rom <= {16'd12368, 16'd30344};
                15'd4038 : data_rom <= {16'd12371, 16'd30342};
                15'd4039 : data_rom <= {16'd12374, 16'd30341};
                15'd4040 : data_rom <= {16'd12377, 16'd30340};
                15'd4041 : data_rom <= {16'd12379, 16'd30339};
                15'd4042 : data_rom <= {16'd12382, 16'd30338};
                15'd4043 : data_rom <= {16'd12385, 16'd30337};
                15'd4044 : data_rom <= {16'd12388, 16'd30335};
                15'd4045 : data_rom <= {16'd12391, 16'd30334};
                15'd4046 : data_rom <= {16'd12394, 16'd30333};
                15'd4047 : data_rom <= {16'd12397, 16'd30332};
                15'd4048 : data_rom <= {16'd12400, 16'd30331};
                15'd4049 : data_rom <= {16'd12403, 16'd30329};
                15'd4050 : data_rom <= {16'd12406, 16'd30328};
                15'd4051 : data_rom <= {16'd12409, 16'd30327};
                15'd4052 : data_rom <= {16'd12411, 16'd30326};
                15'd4053 : data_rom <= {16'd12414, 16'd30325};
                15'd4054 : data_rom <= {16'd12417, 16'd30323};
                15'd4055 : data_rom <= {16'd12420, 16'd30322};
                15'd4056 : data_rom <= {16'd12423, 16'd30321};
                15'd4057 : data_rom <= {16'd12426, 16'd30320};
                15'd4058 : data_rom <= {16'd12429, 16'd30319};
                15'd4059 : data_rom <= {16'd12432, 16'd30317};
                15'd4060 : data_rom <= {16'd12435, 16'd30316};
                15'd4061 : data_rom <= {16'd12438, 16'd30315};
                15'd4062 : data_rom <= {16'd12441, 16'd30314};
                15'd4063 : data_rom <= {16'd12443, 16'd30313};
                15'd4064 : data_rom <= {16'd12446, 16'd30312};
                15'd4065 : data_rom <= {16'd12449, 16'd30310};
                15'd4066 : data_rom <= {16'd12452, 16'd30309};
                15'd4067 : data_rom <= {16'd12455, 16'd30308};
                15'd4068 : data_rom <= {16'd12458, 16'd30307};
                15'd4069 : data_rom <= {16'd12461, 16'd30306};
                15'd4070 : data_rom <= {16'd12464, 16'd30304};
                15'd4071 : data_rom <= {16'd12467, 16'd30303};
                15'd4072 : data_rom <= {16'd12470, 16'd30302};
                15'd4073 : data_rom <= {16'd12472, 16'd30301};
                15'd4074 : data_rom <= {16'd12475, 16'd30300};
                15'd4075 : data_rom <= {16'd12478, 16'd30298};
                15'd4076 : data_rom <= {16'd12481, 16'd30297};
                15'd4077 : data_rom <= {16'd12484, 16'd30296};
                15'd4078 : data_rom <= {16'd12487, 16'd30295};
                15'd4079 : data_rom <= {16'd12490, 16'd30294};
                15'd4080 : data_rom <= {16'd12493, 16'd30292};
                15'd4081 : data_rom <= {16'd12496, 16'd30291};
                15'd4082 : data_rom <= {16'd12499, 16'd30290};
                15'd4083 : data_rom <= {16'd12502, 16'd30289};
                15'd4084 : data_rom <= {16'd12504, 16'd30288};
                15'd4085 : data_rom <= {16'd12507, 16'd30286};
                15'd4086 : data_rom <= {16'd12510, 16'd30285};
                15'd4087 : data_rom <= {16'd12513, 16'd30284};
                15'd4088 : data_rom <= {16'd12516, 16'd30283};
                15'd4089 : data_rom <= {16'd12519, 16'd30282};
                15'd4090 : data_rom <= {16'd12522, 16'd30280};
                15'd4091 : data_rom <= {16'd12525, 16'd30279};
                15'd4092 : data_rom <= {16'd12528, 16'd30278};
                15'd4093 : data_rom <= {16'd12531, 16'd30277};
                15'd4094 : data_rom <= {16'd12533, 16'd30276};
                15'd4095 : data_rom <= {16'd12536, 16'd30274};
                15'd4096 : data_rom <= {16'd12539, 16'd30273};
                15'd4097 : data_rom <= {16'd12542, 16'd30272};
                15'd4098 : data_rom <= {16'd12545, 16'd30271};
                15'd4099 : data_rom <= {16'd12548, 16'd30270};
                15'd4100 : data_rom <= {16'd12551, 16'd30268};
                15'd4101 : data_rom <= {16'd12554, 16'd30267};
                15'd4102 : data_rom <= {16'd12557, 16'd30266};
                15'd4103 : data_rom <= {16'd12560, 16'd30265};
                15'd4104 : data_rom <= {16'd12562, 16'd30264};
                15'd4105 : data_rom <= {16'd12565, 16'd30262};
                15'd4106 : data_rom <= {16'd12568, 16'd30261};
                15'd4107 : data_rom <= {16'd12571, 16'd30260};
                15'd4108 : data_rom <= {16'd12574, 16'd30259};
                15'd4109 : data_rom <= {16'd12577, 16'd30258};
                15'd4110 : data_rom <= {16'd12580, 16'd30256};
                15'd4111 : data_rom <= {16'd12583, 16'd30255};
                15'd4112 : data_rom <= {16'd12586, 16'd30254};
                15'd4113 : data_rom <= {16'd12589, 16'd30253};
                15'd4114 : data_rom <= {16'd12591, 16'd30252};
                15'd4115 : data_rom <= {16'd12594, 16'd30250};
                15'd4116 : data_rom <= {16'd12597, 16'd30249};
                15'd4117 : data_rom <= {16'd12600, 16'd30248};
                15'd4118 : data_rom <= {16'd12603, 16'd30247};
                15'd4119 : data_rom <= {16'd12606, 16'd30245};
                15'd4120 : data_rom <= {16'd12609, 16'd30244};
                15'd4121 : data_rom <= {16'd12612, 16'd30243};
                15'd4122 : data_rom <= {16'd12615, 16'd30242};
                15'd4123 : data_rom <= {16'd12618, 16'd30241};
                15'd4124 : data_rom <= {16'd12620, 16'd30239};
                15'd4125 : data_rom <= {16'd12623, 16'd30238};
                15'd4126 : data_rom <= {16'd12626, 16'd30237};
                15'd4127 : data_rom <= {16'd12629, 16'd30236};
                15'd4128 : data_rom <= {16'd12632, 16'd30235};
                15'd4129 : data_rom <= {16'd12635, 16'd30233};
                15'd4130 : data_rom <= {16'd12638, 16'd30232};
                15'd4131 : data_rom <= {16'd12641, 16'd30231};
                15'd4132 : data_rom <= {16'd12644, 16'd30230};
                15'd4133 : data_rom <= {16'd12647, 16'd30229};
                15'd4134 : data_rom <= {16'd12649, 16'd30227};
                15'd4135 : data_rom <= {16'd12652, 16'd30226};
                15'd4136 : data_rom <= {16'd12655, 16'd30225};
                15'd4137 : data_rom <= {16'd12658, 16'd30224};
                15'd4138 : data_rom <= {16'd12661, 16'd30222};
                15'd4139 : data_rom <= {16'd12664, 16'd30221};
                15'd4140 : data_rom <= {16'd12667, 16'd30220};
                15'd4141 : data_rom <= {16'd12670, 16'd30219};
                15'd4142 : data_rom <= {16'd12673, 16'd30218};
                15'd4143 : data_rom <= {16'd12676, 16'd30216};
                15'd4144 : data_rom <= {16'd12678, 16'd30215};
                15'd4145 : data_rom <= {16'd12681, 16'd30214};
                15'd4146 : data_rom <= {16'd12684, 16'd30213};
                15'd4147 : data_rom <= {16'd12687, 16'd30212};
                15'd4148 : data_rom <= {16'd12690, 16'd30210};
                15'd4149 : data_rom <= {16'd12693, 16'd30209};
                15'd4150 : data_rom <= {16'd12696, 16'd30208};
                15'd4151 : data_rom <= {16'd12699, 16'd30207};
                15'd4152 : data_rom <= {16'd12702, 16'd30205};
                15'd4153 : data_rom <= {16'd12705, 16'd30204};
                15'd4154 : data_rom <= {16'd12707, 16'd30203};
                15'd4155 : data_rom <= {16'd12710, 16'd30202};
                15'd4156 : data_rom <= {16'd12713, 16'd30201};
                15'd4157 : data_rom <= {16'd12716, 16'd30199};
                15'd4158 : data_rom <= {16'd12719, 16'd30198};
                15'd4159 : data_rom <= {16'd12722, 16'd30197};
                15'd4160 : data_rom <= {16'd12725, 16'd30196};
                15'd4161 : data_rom <= {16'd12728, 16'd30194};
                15'd4162 : data_rom <= {16'd12731, 16'd30193};
                15'd4163 : data_rom <= {16'd12733, 16'd30192};
                15'd4164 : data_rom <= {16'd12736, 16'd30191};
                15'd4165 : data_rom <= {16'd12739, 16'd30190};
                15'd4166 : data_rom <= {16'd12742, 16'd30188};
                15'd4167 : data_rom <= {16'd12745, 16'd30187};
                15'd4168 : data_rom <= {16'd12748, 16'd30186};
                15'd4169 : data_rom <= {16'd12751, 16'd30185};
                15'd4170 : data_rom <= {16'd12754, 16'd30183};
                15'd4171 : data_rom <= {16'd12757, 16'd30182};
                15'd4172 : data_rom <= {16'd12760, 16'd30181};
                15'd4173 : data_rom <= {16'd12762, 16'd30180};
                15'd4174 : data_rom <= {16'd12765, 16'd30179};
                15'd4175 : data_rom <= {16'd12768, 16'd30177};
                15'd4176 : data_rom <= {16'd12771, 16'd30176};
                15'd4177 : data_rom <= {16'd12774, 16'd30175};
                15'd4178 : data_rom <= {16'd12777, 16'd30174};
                15'd4179 : data_rom <= {16'd12780, 16'd30172};
                15'd4180 : data_rom <= {16'd12783, 16'd30171};
                15'd4181 : data_rom <= {16'd12786, 16'd30170};
                15'd4182 : data_rom <= {16'd12788, 16'd30169};
                15'd4183 : data_rom <= {16'd12791, 16'd30168};
                15'd4184 : data_rom <= {16'd12794, 16'd30166};
                15'd4185 : data_rom <= {16'd12797, 16'd30165};
                15'd4186 : data_rom <= {16'd12800, 16'd30164};
                15'd4187 : data_rom <= {16'd12803, 16'd30163};
                15'd4188 : data_rom <= {16'd12806, 16'd30161};
                15'd4189 : data_rom <= {16'd12809, 16'd30160};
                15'd4190 : data_rom <= {16'd12812, 16'd30159};
                15'd4191 : data_rom <= {16'd12814, 16'd30158};
                15'd4192 : data_rom <= {16'd12817, 16'd30156};
                15'd4193 : data_rom <= {16'd12820, 16'd30155};
                15'd4194 : data_rom <= {16'd12823, 16'd30154};
                15'd4195 : data_rom <= {16'd12826, 16'd30153};
                15'd4196 : data_rom <= {16'd12829, 16'd30152};
                15'd4197 : data_rom <= {16'd12832, 16'd30150};
                15'd4198 : data_rom <= {16'd12835, 16'd30149};
                15'd4199 : data_rom <= {16'd12838, 16'd30148};
                15'd4200 : data_rom <= {16'd12840, 16'd30147};
                15'd4201 : data_rom <= {16'd12843, 16'd30145};
                15'd4202 : data_rom <= {16'd12846, 16'd30144};
                15'd4203 : data_rom <= {16'd12849, 16'd30143};
                15'd4204 : data_rom <= {16'd12852, 16'd30142};
                15'd4205 : data_rom <= {16'd12855, 16'd30140};
                15'd4206 : data_rom <= {16'd12858, 16'd30139};
                15'd4207 : data_rom <= {16'd12861, 16'd30138};
                15'd4208 : data_rom <= {16'd12864, 16'd30137};
                15'd4209 : data_rom <= {16'd12866, 16'd30136};
                15'd4210 : data_rom <= {16'd12869, 16'd30134};
                15'd4211 : data_rom <= {16'd12872, 16'd30133};
                15'd4212 : data_rom <= {16'd12875, 16'd30132};
                15'd4213 : data_rom <= {16'd12878, 16'd30131};
                15'd4214 : data_rom <= {16'd12881, 16'd30129};
                15'd4215 : data_rom <= {16'd12884, 16'd30128};
                15'd4216 : data_rom <= {16'd12887, 16'd30127};
                15'd4217 : data_rom <= {16'd12890, 16'd30126};
                15'd4218 : data_rom <= {16'd12892, 16'd30124};
                15'd4219 : data_rom <= {16'd12895, 16'd30123};
                15'd4220 : data_rom <= {16'd12898, 16'd30122};
                15'd4221 : data_rom <= {16'd12901, 16'd30121};
                15'd4222 : data_rom <= {16'd12904, 16'd30120};
                15'd4223 : data_rom <= {16'd12907, 16'd30118};
                15'd4224 : data_rom <= {16'd12910, 16'd30117};
                15'd4225 : data_rom <= {16'd12913, 16'd30116};
                15'd4226 : data_rom <= {16'd12916, 16'd30115};
                15'd4227 : data_rom <= {16'd12918, 16'd30113};
                15'd4228 : data_rom <= {16'd12921, 16'd30112};
                15'd4229 : data_rom <= {16'd12924, 16'd30111};
                15'd4230 : data_rom <= {16'd12927, 16'd30110};
                15'd4231 : data_rom <= {16'd12930, 16'd30108};
                15'd4232 : data_rom <= {16'd12933, 16'd30107};
                15'd4233 : data_rom <= {16'd12936, 16'd30106};
                15'd4234 : data_rom <= {16'd12939, 16'd30105};
                15'd4235 : data_rom <= {16'd12942, 16'd30103};
                15'd4236 : data_rom <= {16'd12944, 16'd30102};
                15'd4237 : data_rom <= {16'd12947, 16'd30101};
                15'd4238 : data_rom <= {16'd12950, 16'd30100};
                15'd4239 : data_rom <= {16'd12953, 16'd30098};
                15'd4240 : data_rom <= {16'd12956, 16'd30097};
                15'd4241 : data_rom <= {16'd12959, 16'd30096};
                15'd4242 : data_rom <= {16'd12962, 16'd30095};
                15'd4243 : data_rom <= {16'd12965, 16'd30093};
                15'd4244 : data_rom <= {16'd12968, 16'd30092};
                15'd4245 : data_rom <= {16'd12970, 16'd30091};
                15'd4246 : data_rom <= {16'd12973, 16'd30090};
                15'd4247 : data_rom <= {16'd12976, 16'd30088};
                15'd4248 : data_rom <= {16'd12979, 16'd30087};
                15'd4249 : data_rom <= {16'd12982, 16'd30086};
                15'd4250 : data_rom <= {16'd12985, 16'd30085};
                15'd4251 : data_rom <= {16'd12988, 16'd30084};
                15'd4252 : data_rom <= {16'd12991, 16'd30082};
                15'd4253 : data_rom <= {16'd12994, 16'd30081};
                15'd4254 : data_rom <= {16'd12996, 16'd30080};
                15'd4255 : data_rom <= {16'd12999, 16'd30079};
                15'd4256 : data_rom <= {16'd13002, 16'd30077};
                15'd4257 : data_rom <= {16'd13005, 16'd30076};
                15'd4258 : data_rom <= {16'd13008, 16'd30075};
                15'd4259 : data_rom <= {16'd13011, 16'd30074};
                15'd4260 : data_rom <= {16'd13014, 16'd30072};
                15'd4261 : data_rom <= {16'd13017, 16'd30071};
                15'd4262 : data_rom <= {16'd13019, 16'd30070};
                15'd4263 : data_rom <= {16'd13022, 16'd30069};
                15'd4264 : data_rom <= {16'd13025, 16'd30067};
                15'd4265 : data_rom <= {16'd13028, 16'd30066};
                15'd4266 : data_rom <= {16'd13031, 16'd30065};
                15'd4267 : data_rom <= {16'd13034, 16'd30064};
                15'd4268 : data_rom <= {16'd13037, 16'd30062};
                15'd4269 : data_rom <= {16'd13040, 16'd30061};
                15'd4270 : data_rom <= {16'd13043, 16'd30060};
                15'd4271 : data_rom <= {16'd13045, 16'd30059};
                15'd4272 : data_rom <= {16'd13048, 16'd30057};
                15'd4273 : data_rom <= {16'd13051, 16'd30056};
                15'd4274 : data_rom <= {16'd13054, 16'd30055};
                15'd4275 : data_rom <= {16'd13057, 16'd30054};
                15'd4276 : data_rom <= {16'd13060, 16'd30052};
                15'd4277 : data_rom <= {16'd13063, 16'd30051};
                15'd4278 : data_rom <= {16'd13066, 16'd30050};
                15'd4279 : data_rom <= {16'd13068, 16'd30049};
                15'd4280 : data_rom <= {16'd13071, 16'd30047};
                15'd4281 : data_rom <= {16'd13074, 16'd30046};
                15'd4282 : data_rom <= {16'd13077, 16'd30045};
                15'd4283 : data_rom <= {16'd13080, 16'd30044};
                15'd4284 : data_rom <= {16'd13083, 16'd30042};
                15'd4285 : data_rom <= {16'd13086, 16'd30041};
                15'd4286 : data_rom <= {16'd13089, 16'd30040};
                15'd4287 : data_rom <= {16'd13091, 16'd30038};
                15'd4288 : data_rom <= {16'd13094, 16'd30037};
                15'd4289 : data_rom <= {16'd13097, 16'd30036};
                15'd4290 : data_rom <= {16'd13100, 16'd30035};
                15'd4291 : data_rom <= {16'd13103, 16'd30033};
                15'd4292 : data_rom <= {16'd13106, 16'd30032};
                15'd4293 : data_rom <= {16'd13109, 16'd30031};
                15'd4294 : data_rom <= {16'd13112, 16'd30030};
                15'd4295 : data_rom <= {16'd13115, 16'd30028};
                15'd4296 : data_rom <= {16'd13117, 16'd30027};
                15'd4297 : data_rom <= {16'd13120, 16'd30026};
                15'd4298 : data_rom <= {16'd13123, 16'd30025};
                15'd4299 : data_rom <= {16'd13126, 16'd30023};
                15'd4300 : data_rom <= {16'd13129, 16'd30022};
                15'd4301 : data_rom <= {16'd13132, 16'd30021};
                15'd4302 : data_rom <= {16'd13135, 16'd30020};
                15'd4303 : data_rom <= {16'd13138, 16'd30018};
                15'd4304 : data_rom <= {16'd13140, 16'd30017};
                15'd4305 : data_rom <= {16'd13143, 16'd30016};
                15'd4306 : data_rom <= {16'd13146, 16'd30015};
                15'd4307 : data_rom <= {16'd13149, 16'd30013};
                15'd4308 : data_rom <= {16'd13152, 16'd30012};
                15'd4309 : data_rom <= {16'd13155, 16'd30011};
                15'd4310 : data_rom <= {16'd13158, 16'd30010};
                15'd4311 : data_rom <= {16'd13161, 16'd30008};
                15'd4312 : data_rom <= {16'd13163, 16'd30007};
                15'd4313 : data_rom <= {16'd13166, 16'd30006};
                15'd4314 : data_rom <= {16'd13169, 16'd30005};
                15'd4315 : data_rom <= {16'd13172, 16'd30003};
                15'd4316 : data_rom <= {16'd13175, 16'd30002};
                15'd4317 : data_rom <= {16'd13178, 16'd30001};
                15'd4318 : data_rom <= {16'd13181, 16'd29999};
                15'd4319 : data_rom <= {16'd13184, 16'd29998};
                15'd4320 : data_rom <= {16'd13186, 16'd29997};
                15'd4321 : data_rom <= {16'd13189, 16'd29996};
                15'd4322 : data_rom <= {16'd13192, 16'd29994};
                15'd4323 : data_rom <= {16'd13195, 16'd29993};
                15'd4324 : data_rom <= {16'd13198, 16'd29992};
                15'd4325 : data_rom <= {16'd13201, 16'd29991};
                15'd4326 : data_rom <= {16'd13204, 16'd29989};
                15'd4327 : data_rom <= {16'd13207, 16'd29988};
                15'd4328 : data_rom <= {16'd13209, 16'd29987};
                15'd4329 : data_rom <= {16'd13212, 16'd29986};
                15'd4330 : data_rom <= {16'd13215, 16'd29984};
                15'd4331 : data_rom <= {16'd13218, 16'd29983};
                15'd4332 : data_rom <= {16'd13221, 16'd29982};
                15'd4333 : data_rom <= {16'd13224, 16'd29980};
                15'd4334 : data_rom <= {16'd13227, 16'd29979};
                15'd4335 : data_rom <= {16'd13230, 16'd29978};
                15'd4336 : data_rom <= {16'd13232, 16'd29977};
                15'd4337 : data_rom <= {16'd13235, 16'd29975};
                15'd4338 : data_rom <= {16'd13238, 16'd29974};
                15'd4339 : data_rom <= {16'd13241, 16'd29973};
                15'd4340 : data_rom <= {16'd13244, 16'd29972};
                15'd4341 : data_rom <= {16'd13247, 16'd29970};
                15'd4342 : data_rom <= {16'd13250, 16'd29969};
                15'd4343 : data_rom <= {16'd13253, 16'd29968};
                15'd4344 : data_rom <= {16'd13255, 16'd29967};
                15'd4345 : data_rom <= {16'd13258, 16'd29965};
                15'd4346 : data_rom <= {16'd13261, 16'd29964};
                15'd4347 : data_rom <= {16'd13264, 16'd29963};
                15'd4348 : data_rom <= {16'd13267, 16'd29961};
                15'd4349 : data_rom <= {16'd13270, 16'd29960};
                15'd4350 : data_rom <= {16'd13273, 16'd29959};
                15'd4351 : data_rom <= {16'd13276, 16'd29958};
                15'd4352 : data_rom <= {16'd13278, 16'd29956};
                15'd4353 : data_rom <= {16'd13281, 16'd29955};
                15'd4354 : data_rom <= {16'd13284, 16'd29954};
                15'd4355 : data_rom <= {16'd13287, 16'd29953};
                15'd4356 : data_rom <= {16'd13290, 16'd29951};
                15'd4357 : data_rom <= {16'd13293, 16'd29950};
                15'd4358 : data_rom <= {16'd13296, 16'd29949};
                15'd4359 : data_rom <= {16'd13299, 16'd29947};
                15'd4360 : data_rom <= {16'd13301, 16'd29946};
                15'd4361 : data_rom <= {16'd13304, 16'd29945};
                15'd4362 : data_rom <= {16'd13307, 16'd29944};
                15'd4363 : data_rom <= {16'd13310, 16'd29942};
                15'd4364 : data_rom <= {16'd13313, 16'd29941};
                15'd4365 : data_rom <= {16'd13316, 16'd29940};
                15'd4366 : data_rom <= {16'd13319, 16'd29938};
                15'd4367 : data_rom <= {16'd13322, 16'd29937};
                15'd4368 : data_rom <= {16'd13324, 16'd29936};
                15'd4369 : data_rom <= {16'd13327, 16'd29935};
                15'd4370 : data_rom <= {16'd13330, 16'd29933};
                15'd4371 : data_rom <= {16'd13333, 16'd29932};
                15'd4372 : data_rom <= {16'd13336, 16'd29931};
                15'd4373 : data_rom <= {16'd13339, 16'd29930};
                15'd4374 : data_rom <= {16'd13342, 16'd29928};
                15'd4375 : data_rom <= {16'd13344, 16'd29927};
                15'd4376 : data_rom <= {16'd13347, 16'd29926};
                15'd4377 : data_rom <= {16'd13350, 16'd29924};
                15'd4378 : data_rom <= {16'd13353, 16'd29923};
                15'd4379 : data_rom <= {16'd13356, 16'd29922};
                15'd4380 : data_rom <= {16'd13359, 16'd29921};
                15'd4381 : data_rom <= {16'd13362, 16'd29919};
                15'd4382 : data_rom <= {16'd13365, 16'd29918};
                15'd4383 : data_rom <= {16'd13367, 16'd29917};
                15'd4384 : data_rom <= {16'd13370, 16'd29915};
                15'd4385 : data_rom <= {16'd13373, 16'd29914};
                15'd4386 : data_rom <= {16'd13376, 16'd29913};
                15'd4387 : data_rom <= {16'd13379, 16'd29912};
                15'd4388 : data_rom <= {16'd13382, 16'd29910};
                15'd4389 : data_rom <= {16'd13385, 16'd29909};
                15'd4390 : data_rom <= {16'd13387, 16'd29908};
                15'd4391 : data_rom <= {16'd13390, 16'd29906};
                15'd4392 : data_rom <= {16'd13393, 16'd29905};
                15'd4393 : data_rom <= {16'd13396, 16'd29904};
                15'd4394 : data_rom <= {16'd13399, 16'd29903};
                15'd4395 : data_rom <= {16'd13402, 16'd29901};
                15'd4396 : data_rom <= {16'd13405, 16'd29900};
                15'd4397 : data_rom <= {16'd13408, 16'd29899};
                15'd4398 : data_rom <= {16'd13410, 16'd29897};
                15'd4399 : data_rom <= {16'd13413, 16'd29896};
                15'd4400 : data_rom <= {16'd13416, 16'd29895};
                15'd4401 : data_rom <= {16'd13419, 16'd29894};
                15'd4402 : data_rom <= {16'd13422, 16'd29892};
                15'd4403 : data_rom <= {16'd13425, 16'd29891};
                15'd4404 : data_rom <= {16'd13428, 16'd29890};
                15'd4405 : data_rom <= {16'd13430, 16'd29888};
                15'd4406 : data_rom <= {16'd13433, 16'd29887};
                15'd4407 : data_rom <= {16'd13436, 16'd29886};
                15'd4408 : data_rom <= {16'd13439, 16'd29885};
                15'd4409 : data_rom <= {16'd13442, 16'd29883};
                15'd4410 : data_rom <= {16'd13445, 16'd29882};
                15'd4411 : data_rom <= {16'd13448, 16'd29881};
                15'd4412 : data_rom <= {16'd13451, 16'd29879};
                15'd4413 : data_rom <= {16'd13453, 16'd29878};
                15'd4414 : data_rom <= {16'd13456, 16'd29877};
                15'd4415 : data_rom <= {16'd13459, 16'd29876};
                15'd4416 : data_rom <= {16'd13462, 16'd29874};
                15'd4417 : data_rom <= {16'd13465, 16'd29873};
                15'd4418 : data_rom <= {16'd13468, 16'd29872};
                15'd4419 : data_rom <= {16'd13471, 16'd29870};
                15'd4420 : data_rom <= {16'd13473, 16'd29869};
                15'd4421 : data_rom <= {16'd13476, 16'd29868};
                15'd4422 : data_rom <= {16'd13479, 16'd29867};
                15'd4423 : data_rom <= {16'd13482, 16'd29865};
                15'd4424 : data_rom <= {16'd13485, 16'd29864};
                15'd4425 : data_rom <= {16'd13488, 16'd29863};
                15'd4426 : data_rom <= {16'd13491, 16'd29861};
                15'd4427 : data_rom <= {16'd13493, 16'd29860};
                15'd4428 : data_rom <= {16'd13496, 16'd29859};
                15'd4429 : data_rom <= {16'd13499, 16'd29857};
                15'd4430 : data_rom <= {16'd13502, 16'd29856};
                15'd4431 : data_rom <= {16'd13505, 16'd29855};
                15'd4432 : data_rom <= {16'd13508, 16'd29854};
                15'd4433 : data_rom <= {16'd13511, 16'd29852};
                15'd4434 : data_rom <= {16'd13514, 16'd29851};
                15'd4435 : data_rom <= {16'd13516, 16'd29850};
                15'd4436 : data_rom <= {16'd13519, 16'd29848};
                15'd4437 : data_rom <= {16'd13522, 16'd29847};
                15'd4438 : data_rom <= {16'd13525, 16'd29846};
                15'd4439 : data_rom <= {16'd13528, 16'd29845};
                15'd4440 : data_rom <= {16'd13531, 16'd29843};
                15'd4441 : data_rom <= {16'd13534, 16'd29842};
                15'd4442 : data_rom <= {16'd13536, 16'd29841};
                15'd4443 : data_rom <= {16'd13539, 16'd29839};
                15'd4444 : data_rom <= {16'd13542, 16'd29838};
                15'd4445 : data_rom <= {16'd13545, 16'd29837};
                15'd4446 : data_rom <= {16'd13548, 16'd29835};
                15'd4447 : data_rom <= {16'd13551, 16'd29834};
                15'd4448 : data_rom <= {16'd13554, 16'd29833};
                15'd4449 : data_rom <= {16'd13556, 16'd29832};
                15'd4450 : data_rom <= {16'd13559, 16'd29830};
                15'd4451 : data_rom <= {16'd13562, 16'd29829};
                15'd4452 : data_rom <= {16'd13565, 16'd29828};
                15'd4453 : data_rom <= {16'd13568, 16'd29826};
                15'd4454 : data_rom <= {16'd13571, 16'd29825};
                15'd4455 : data_rom <= {16'd13574, 16'd29824};
                15'd4456 : data_rom <= {16'd13576, 16'd29822};
                15'd4457 : data_rom <= {16'd13579, 16'd29821};
                15'd4458 : data_rom <= {16'd13582, 16'd29820};
                15'd4459 : data_rom <= {16'd13585, 16'd29819};
                15'd4460 : data_rom <= {16'd13588, 16'd29817};
                15'd4461 : data_rom <= {16'd13591, 16'd29816};
                15'd4462 : data_rom <= {16'd13594, 16'd29815};
                15'd4463 : data_rom <= {16'd13596, 16'd29813};
                15'd4464 : data_rom <= {16'd13599, 16'd29812};
                15'd4465 : data_rom <= {16'd13602, 16'd29811};
                15'd4466 : data_rom <= {16'd13605, 16'd29809};
                15'd4467 : data_rom <= {16'd13608, 16'd29808};
                15'd4468 : data_rom <= {16'd13611, 16'd29807};
                15'd4469 : data_rom <= {16'd13614, 16'd29805};
                15'd4470 : data_rom <= {16'd13616, 16'd29804};
                15'd4471 : data_rom <= {16'd13619, 16'd29803};
                15'd4472 : data_rom <= {16'd13622, 16'd29802};
                15'd4473 : data_rom <= {16'd13625, 16'd29800};
                15'd4474 : data_rom <= {16'd13628, 16'd29799};
                15'd4475 : data_rom <= {16'd13631, 16'd29798};
                15'd4476 : data_rom <= {16'd13634, 16'd29796};
                15'd4477 : data_rom <= {16'd13636, 16'd29795};
                15'd4478 : data_rom <= {16'd13639, 16'd29794};
                15'd4479 : data_rom <= {16'd13642, 16'd29792};
                15'd4480 : data_rom <= {16'd13645, 16'd29791};
                15'd4481 : data_rom <= {16'd13648, 16'd29790};
                15'd4482 : data_rom <= {16'd13651, 16'd29789};
                15'd4483 : data_rom <= {16'd13654, 16'd29787};
                15'd4484 : data_rom <= {16'd13656, 16'd29786};
                15'd4485 : data_rom <= {16'd13659, 16'd29785};
                15'd4486 : data_rom <= {16'd13662, 16'd29783};
                15'd4487 : data_rom <= {16'd13665, 16'd29782};
                15'd4488 : data_rom <= {16'd13668, 16'd29781};
                15'd4489 : data_rom <= {16'd13671, 16'd29779};
                15'd4490 : data_rom <= {16'd13674, 16'd29778};
                15'd4491 : data_rom <= {16'd13676, 16'd29777};
                15'd4492 : data_rom <= {16'd13679, 16'd29775};
                15'd4493 : data_rom <= {16'd13682, 16'd29774};
                15'd4494 : data_rom <= {16'd13685, 16'd29773};
                15'd4495 : data_rom <= {16'd13688, 16'd29771};
                15'd4496 : data_rom <= {16'd13691, 16'd29770};
                15'd4497 : data_rom <= {16'd13694, 16'd29769};
                15'd4498 : data_rom <= {16'd13696, 16'd29768};
                15'd4499 : data_rom <= {16'd13699, 16'd29766};
                15'd4500 : data_rom <= {16'd13702, 16'd29765};
                15'd4501 : data_rom <= {16'd13705, 16'd29764};
                15'd4502 : data_rom <= {16'd13708, 16'd29762};
                15'd4503 : data_rom <= {16'd13711, 16'd29761};
                15'd4504 : data_rom <= {16'd13714, 16'd29760};
                15'd4505 : data_rom <= {16'd13716, 16'd29758};
                15'd4506 : data_rom <= {16'd13719, 16'd29757};
                15'd4507 : data_rom <= {16'd13722, 16'd29756};
                15'd4508 : data_rom <= {16'd13725, 16'd29754};
                15'd4509 : data_rom <= {16'd13728, 16'd29753};
                15'd4510 : data_rom <= {16'd13731, 16'd29752};
                15'd4511 : data_rom <= {16'd13734, 16'd29750};
                15'd4512 : data_rom <= {16'd13736, 16'd29749};
                15'd4513 : data_rom <= {16'd13739, 16'd29748};
                15'd4514 : data_rom <= {16'd13742, 16'd29746};
                15'd4515 : data_rom <= {16'd13745, 16'd29745};
                15'd4516 : data_rom <= {16'd13748, 16'd29744};
                15'd4517 : data_rom <= {16'd13751, 16'd29743};
                15'd4518 : data_rom <= {16'd13753, 16'd29741};
                15'd4519 : data_rom <= {16'd13756, 16'd29740};
                15'd4520 : data_rom <= {16'd13759, 16'd29739};
                15'd4521 : data_rom <= {16'd13762, 16'd29737};
                15'd4522 : data_rom <= {16'd13765, 16'd29736};
                15'd4523 : data_rom <= {16'd13768, 16'd29735};
                15'd4524 : data_rom <= {16'd13771, 16'd29733};
                15'd4525 : data_rom <= {16'd13773, 16'd29732};
                15'd4526 : data_rom <= {16'd13776, 16'd29731};
                15'd4527 : data_rom <= {16'd13779, 16'd29729};
                15'd4528 : data_rom <= {16'd13782, 16'd29728};
                15'd4529 : data_rom <= {16'd13785, 16'd29727};
                15'd4530 : data_rom <= {16'd13788, 16'd29725};
                15'd4531 : data_rom <= {16'd13791, 16'd29724};
                15'd4532 : data_rom <= {16'd13793, 16'd29723};
                15'd4533 : data_rom <= {16'd13796, 16'd29721};
                15'd4534 : data_rom <= {16'd13799, 16'd29720};
                15'd4535 : data_rom <= {16'd13802, 16'd29719};
                15'd4536 : data_rom <= {16'd13805, 16'd29717};
                15'd4537 : data_rom <= {16'd13808, 16'd29716};
                15'd4538 : data_rom <= {16'd13811, 16'd29715};
                15'd4539 : data_rom <= {16'd13813, 16'd29713};
                15'd4540 : data_rom <= {16'd13816, 16'd29712};
                15'd4541 : data_rom <= {16'd13819, 16'd29711};
                15'd4542 : data_rom <= {16'd13822, 16'd29709};
                15'd4543 : data_rom <= {16'd13825, 16'd29708};
                15'd4544 : data_rom <= {16'd13828, 16'd29707};
                15'd4545 : data_rom <= {16'd13830, 16'd29706};
                15'd4546 : data_rom <= {16'd13833, 16'd29704};
                15'd4547 : data_rom <= {16'd13836, 16'd29703};
                15'd4548 : data_rom <= {16'd13839, 16'd29702};
                15'd4549 : data_rom <= {16'd13842, 16'd29700};
                15'd4550 : data_rom <= {16'd13845, 16'd29699};
                15'd4551 : data_rom <= {16'd13848, 16'd29698};
                15'd4552 : data_rom <= {16'd13850, 16'd29696};
                15'd4553 : data_rom <= {16'd13853, 16'd29695};
                15'd4554 : data_rom <= {16'd13856, 16'd29694};
                15'd4555 : data_rom <= {16'd13859, 16'd29692};
                15'd4556 : data_rom <= {16'd13862, 16'd29691};
                15'd4557 : data_rom <= {16'd13865, 16'd29690};
                15'd4558 : data_rom <= {16'd13867, 16'd29688};
                15'd4559 : data_rom <= {16'd13870, 16'd29687};
                15'd4560 : data_rom <= {16'd13873, 16'd29686};
                15'd4561 : data_rom <= {16'd13876, 16'd29684};
                15'd4562 : data_rom <= {16'd13879, 16'd29683};
                15'd4563 : data_rom <= {16'd13882, 16'd29682};
                15'd4564 : data_rom <= {16'd13885, 16'd29680};
                15'd4565 : data_rom <= {16'd13887, 16'd29679};
                15'd4566 : data_rom <= {16'd13890, 16'd29678};
                15'd4567 : data_rom <= {16'd13893, 16'd29676};
                15'd4568 : data_rom <= {16'd13896, 16'd29675};
                15'd4569 : data_rom <= {16'd13899, 16'd29674};
                15'd4570 : data_rom <= {16'd13902, 16'd29672};
                15'd4571 : data_rom <= {16'd13904, 16'd29671};
                15'd4572 : data_rom <= {16'd13907, 16'd29670};
                15'd4573 : data_rom <= {16'd13910, 16'd29668};
                15'd4574 : data_rom <= {16'd13913, 16'd29667};
                15'd4575 : data_rom <= {16'd13916, 16'd29666};
                15'd4576 : data_rom <= {16'd13919, 16'd29664};
                15'd4577 : data_rom <= {16'd13922, 16'd29663};
                15'd4578 : data_rom <= {16'd13924, 16'd29662};
                15'd4579 : data_rom <= {16'd13927, 16'd29660};
                15'd4580 : data_rom <= {16'd13930, 16'd29659};
                15'd4581 : data_rom <= {16'd13933, 16'd29658};
                15'd4582 : data_rom <= {16'd13936, 16'd29656};
                15'd4583 : data_rom <= {16'd13939, 16'd29655};
                15'd4584 : data_rom <= {16'd13941, 16'd29654};
                15'd4585 : data_rom <= {16'd13944, 16'd29652};
                15'd4586 : data_rom <= {16'd13947, 16'd29651};
                15'd4587 : data_rom <= {16'd13950, 16'd29650};
                15'd4588 : data_rom <= {16'd13953, 16'd29648};
                15'd4589 : data_rom <= {16'd13956, 16'd29647};
                15'd4590 : data_rom <= {16'd13958, 16'd29646};
                15'd4591 : data_rom <= {16'd13961, 16'd29644};
                15'd4592 : data_rom <= {16'd13964, 16'd29643};
                15'd4593 : data_rom <= {16'd13967, 16'd29642};
                15'd4594 : data_rom <= {16'd13970, 16'd29640};
                15'd4595 : data_rom <= {16'd13973, 16'd29639};
                15'd4596 : data_rom <= {16'd13976, 16'd29638};
                15'd4597 : data_rom <= {16'd13978, 16'd29636};
                15'd4598 : data_rom <= {16'd13981, 16'd29635};
                15'd4599 : data_rom <= {16'd13984, 16'd29634};
                15'd4600 : data_rom <= {16'd13987, 16'd29632};
                15'd4601 : data_rom <= {16'd13990, 16'd29631};
                15'd4602 : data_rom <= {16'd13993, 16'd29629};
                15'd4603 : data_rom <= {16'd13995, 16'd29628};
                15'd4604 : data_rom <= {16'd13998, 16'd29627};
                15'd4605 : data_rom <= {16'd14001, 16'd29625};
                15'd4606 : data_rom <= {16'd14004, 16'd29624};
                15'd4607 : data_rom <= {16'd14007, 16'd29623};
                15'd4608 : data_rom <= {16'd14010, 16'd29621};
                15'd4609 : data_rom <= {16'd14012, 16'd29620};
                15'd4610 : data_rom <= {16'd14015, 16'd29619};
                15'd4611 : data_rom <= {16'd14018, 16'd29617};
                15'd4612 : data_rom <= {16'd14021, 16'd29616};
                15'd4613 : data_rom <= {16'd14024, 16'd29615};
                15'd4614 : data_rom <= {16'd14027, 16'd29613};
                15'd4615 : data_rom <= {16'd14029, 16'd29612};
                15'd4616 : data_rom <= {16'd14032, 16'd29611};
                15'd4617 : data_rom <= {16'd14035, 16'd29609};
                15'd4618 : data_rom <= {16'd14038, 16'd29608};
                15'd4619 : data_rom <= {16'd14041, 16'd29607};
                15'd4620 : data_rom <= {16'd14044, 16'd29605};
                15'd4621 : data_rom <= {16'd14047, 16'd29604};
                15'd4622 : data_rom <= {16'd14049, 16'd29603};
                15'd4623 : data_rom <= {16'd14052, 16'd29601};
                15'd4624 : data_rom <= {16'd14055, 16'd29600};
                15'd4625 : data_rom <= {16'd14058, 16'd29599};
                15'd4626 : data_rom <= {16'd14061, 16'd29597};
                15'd4627 : data_rom <= {16'd14064, 16'd29596};
                15'd4628 : data_rom <= {16'd14066, 16'd29595};
                15'd4629 : data_rom <= {16'd14069, 16'd29593};
                15'd4630 : data_rom <= {16'd14072, 16'd29592};
                15'd4631 : data_rom <= {16'd14075, 16'd29590};
                15'd4632 : data_rom <= {16'd14078, 16'd29589};
                15'd4633 : data_rom <= {16'd14081, 16'd29588};
                15'd4634 : data_rom <= {16'd14083, 16'd29586};
                15'd4635 : data_rom <= {16'd14086, 16'd29585};
                15'd4636 : data_rom <= {16'd14089, 16'd29584};
                15'd4637 : data_rom <= {16'd14092, 16'd29582};
                15'd4638 : data_rom <= {16'd14095, 16'd29581};
                15'd4639 : data_rom <= {16'd14098, 16'd29580};
                15'd4640 : data_rom <= {16'd14100, 16'd29578};
                15'd4641 : data_rom <= {16'd14103, 16'd29577};
                15'd4642 : data_rom <= {16'd14106, 16'd29576};
                15'd4643 : data_rom <= {16'd14109, 16'd29574};
                15'd4644 : data_rom <= {16'd14112, 16'd29573};
                15'd4645 : data_rom <= {16'd14115, 16'd29572};
                15'd4646 : data_rom <= {16'd14117, 16'd29570};
                15'd4647 : data_rom <= {16'd14120, 16'd29569};
                15'd4648 : data_rom <= {16'd14123, 16'd29567};
                15'd4649 : data_rom <= {16'd14126, 16'd29566};
                15'd4650 : data_rom <= {16'd14129, 16'd29565};
                15'd4651 : data_rom <= {16'd14132, 16'd29563};
                15'd4652 : data_rom <= {16'd14134, 16'd29562};
                15'd4653 : data_rom <= {16'd14137, 16'd29561};
                15'd4654 : data_rom <= {16'd14140, 16'd29559};
                15'd4655 : data_rom <= {16'd14143, 16'd29558};
                15'd4656 : data_rom <= {16'd14146, 16'd29557};
                15'd4657 : data_rom <= {16'd14149, 16'd29555};
                15'd4658 : data_rom <= {16'd14151, 16'd29554};
                15'd4659 : data_rom <= {16'd14154, 16'd29553};
                15'd4660 : data_rom <= {16'd14157, 16'd29551};
                15'd4661 : data_rom <= {16'd14160, 16'd29550};
                15'd4662 : data_rom <= {16'd14163, 16'd29548};
                15'd4663 : data_rom <= {16'd14166, 16'd29547};
                15'd4664 : data_rom <= {16'd14168, 16'd29546};
                15'd4665 : data_rom <= {16'd14171, 16'd29544};
                15'd4666 : data_rom <= {16'd14174, 16'd29543};
                15'd4667 : data_rom <= {16'd14177, 16'd29542};
                15'd4668 : data_rom <= {16'd14180, 16'd29540};
                15'd4669 : data_rom <= {16'd14183, 16'd29539};
                15'd4670 : data_rom <= {16'd14185, 16'd29538};
                15'd4671 : data_rom <= {16'd14188, 16'd29536};
                15'd4672 : data_rom <= {16'd14191, 16'd29535};
                15'd4673 : data_rom <= {16'd14194, 16'd29534};
                15'd4674 : data_rom <= {16'd14197, 16'd29532};
                15'd4675 : data_rom <= {16'd14200, 16'd29531};
                15'd4676 : data_rom <= {16'd14202, 16'd29529};
                15'd4677 : data_rom <= {16'd14205, 16'd29528};
                15'd4678 : data_rom <= {16'd14208, 16'd29527};
                15'd4679 : data_rom <= {16'd14211, 16'd29525};
                15'd4680 : data_rom <= {16'd14214, 16'd29524};
                15'd4681 : data_rom <= {16'd14217, 16'd29523};
                15'd4682 : data_rom <= {16'd14219, 16'd29521};
                15'd4683 : data_rom <= {16'd14222, 16'd29520};
                15'd4684 : data_rom <= {16'd14225, 16'd29519};
                15'd4685 : data_rom <= {16'd14228, 16'd29517};
                15'd4686 : data_rom <= {16'd14231, 16'd29516};
                15'd4687 : data_rom <= {16'd14234, 16'd29514};
                15'd4688 : data_rom <= {16'd14236, 16'd29513};
                15'd4689 : data_rom <= {16'd14239, 16'd29512};
                15'd4690 : data_rom <= {16'd14242, 16'd29510};
                15'd4691 : data_rom <= {16'd14245, 16'd29509};
                15'd4692 : data_rom <= {16'd14248, 16'd29508};
                15'd4693 : data_rom <= {16'd14251, 16'd29506};
                15'd4694 : data_rom <= {16'd14253, 16'd29505};
                15'd4695 : data_rom <= {16'd14256, 16'd29504};
                15'd4696 : data_rom <= {16'd14259, 16'd29502};
                15'd4697 : data_rom <= {16'd14262, 16'd29501};
                15'd4698 : data_rom <= {16'd14265, 16'd29499};
                15'd4699 : data_rom <= {16'd14268, 16'd29498};
                15'd4700 : data_rom <= {16'd14270, 16'd29497};
                15'd4701 : data_rom <= {16'd14273, 16'd29495};
                15'd4702 : data_rom <= {16'd14276, 16'd29494};
                15'd4703 : data_rom <= {16'd14279, 16'd29493};
                15'd4704 : data_rom <= {16'd14282, 16'd29491};
                15'd4705 : data_rom <= {16'd14284, 16'd29490};
                15'd4706 : data_rom <= {16'd14287, 16'd29488};
                15'd4707 : data_rom <= {16'd14290, 16'd29487};
                15'd4708 : data_rom <= {16'd14293, 16'd29486};
                15'd4709 : data_rom <= {16'd14296, 16'd29484};
                15'd4710 : data_rom <= {16'd14299, 16'd29483};
                15'd4711 : data_rom <= {16'd14301, 16'd29482};
                15'd4712 : data_rom <= {16'd14304, 16'd29480};
                15'd4713 : data_rom <= {16'd14307, 16'd29479};
                15'd4714 : data_rom <= {16'd14310, 16'd29478};
                15'd4715 : data_rom <= {16'd14313, 16'd29476};
                15'd4716 : data_rom <= {16'd14316, 16'd29475};
                15'd4717 : data_rom <= {16'd14318, 16'd29473};
                15'd4718 : data_rom <= {16'd14321, 16'd29472};
                15'd4719 : data_rom <= {16'd14324, 16'd29471};
                15'd4720 : data_rom <= {16'd14327, 16'd29469};
                15'd4721 : data_rom <= {16'd14330, 16'd29468};
                15'd4722 : data_rom <= {16'd14333, 16'd29467};
                15'd4723 : data_rom <= {16'd14335, 16'd29465};
                15'd4724 : data_rom <= {16'd14338, 16'd29464};
                15'd4725 : data_rom <= {16'd14341, 16'd29462};
                15'd4726 : data_rom <= {16'd14344, 16'd29461};
                15'd4727 : data_rom <= {16'd14347, 16'd29460};
                15'd4728 : data_rom <= {16'd14349, 16'd29458};
                15'd4729 : data_rom <= {16'd14352, 16'd29457};
                15'd4730 : data_rom <= {16'd14355, 16'd29456};
                15'd4731 : data_rom <= {16'd14358, 16'd29454};
                15'd4732 : data_rom <= {16'd14361, 16'd29453};
                15'd4733 : data_rom <= {16'd14364, 16'd29451};
                15'd4734 : data_rom <= {16'd14366, 16'd29450};
                15'd4735 : data_rom <= {16'd14369, 16'd29449};
                15'd4736 : data_rom <= {16'd14372, 16'd29447};
                15'd4737 : data_rom <= {16'd14375, 16'd29446};
                15'd4738 : data_rom <= {16'd14378, 16'd29445};
                15'd4739 : data_rom <= {16'd14381, 16'd29443};
                15'd4740 : data_rom <= {16'd14383, 16'd29442};
                15'd4741 : data_rom <= {16'd14386, 16'd29440};
                15'd4742 : data_rom <= {16'd14389, 16'd29439};
                15'd4743 : data_rom <= {16'd14392, 16'd29438};
                15'd4744 : data_rom <= {16'd14395, 16'd29436};
                15'd4745 : data_rom <= {16'd14397, 16'd29435};
                15'd4746 : data_rom <= {16'd14400, 16'd29433};
                15'd4747 : data_rom <= {16'd14403, 16'd29432};
                15'd4748 : data_rom <= {16'd14406, 16'd29431};
                15'd4749 : data_rom <= {16'd14409, 16'd29429};
                15'd4750 : data_rom <= {16'd14412, 16'd29428};
                15'd4751 : data_rom <= {16'd14414, 16'd29427};
                15'd4752 : data_rom <= {16'd14417, 16'd29425};
                15'd4753 : data_rom <= {16'd14420, 16'd29424};
                15'd4754 : data_rom <= {16'd14423, 16'd29422};
                15'd4755 : data_rom <= {16'd14426, 16'd29421};
                15'd4756 : data_rom <= {16'd14429, 16'd29420};
                15'd4757 : data_rom <= {16'd14431, 16'd29418};
                15'd4758 : data_rom <= {16'd14434, 16'd29417};
                15'd4759 : data_rom <= {16'd14437, 16'd29416};
                15'd4760 : data_rom <= {16'd14440, 16'd29414};
                15'd4761 : data_rom <= {16'd14443, 16'd29413};
                15'd4762 : data_rom <= {16'd14445, 16'd29411};
                15'd4763 : data_rom <= {16'd14448, 16'd29410};
                15'd4764 : data_rom <= {16'd14451, 16'd29409};
                15'd4765 : data_rom <= {16'd14454, 16'd29407};
                15'd4766 : data_rom <= {16'd14457, 16'd29406};
                15'd4767 : data_rom <= {16'd14460, 16'd29404};
                15'd4768 : data_rom <= {16'd14462, 16'd29403};
                15'd4769 : data_rom <= {16'd14465, 16'd29402};
                15'd4770 : data_rom <= {16'd14468, 16'd29400};
                15'd4771 : data_rom <= {16'd14471, 16'd29399};
                15'd4772 : data_rom <= {16'd14474, 16'd29397};
                15'd4773 : data_rom <= {16'd14476, 16'd29396};
                15'd4774 : data_rom <= {16'd14479, 16'd29395};
                15'd4775 : data_rom <= {16'd14482, 16'd29393};
                15'd4776 : data_rom <= {16'd14485, 16'd29392};
                15'd4777 : data_rom <= {16'd14488, 16'd29391};
                15'd4778 : data_rom <= {16'd14491, 16'd29389};
                15'd4779 : data_rom <= {16'd14493, 16'd29388};
                15'd4780 : data_rom <= {16'd14496, 16'd29386};
                15'd4781 : data_rom <= {16'd14499, 16'd29385};
                15'd4782 : data_rom <= {16'd14502, 16'd29384};
                15'd4783 : data_rom <= {16'd14505, 16'd29382};
                15'd4784 : data_rom <= {16'd14507, 16'd29381};
                15'd4785 : data_rom <= {16'd14510, 16'd29379};
                15'd4786 : data_rom <= {16'd14513, 16'd29378};
                15'd4787 : data_rom <= {16'd14516, 16'd29377};
                15'd4788 : data_rom <= {16'd14519, 16'd29375};
                15'd4789 : data_rom <= {16'd14522, 16'd29374};
                15'd4790 : data_rom <= {16'd14524, 16'd29372};
                15'd4791 : data_rom <= {16'd14527, 16'd29371};
                15'd4792 : data_rom <= {16'd14530, 16'd29370};
                15'd4793 : data_rom <= {16'd14533, 16'd29368};
                15'd4794 : data_rom <= {16'd14536, 16'd29367};
                15'd4795 : data_rom <= {16'd14538, 16'd29366};
                15'd4796 : data_rom <= {16'd14541, 16'd29364};
                15'd4797 : data_rom <= {16'd14544, 16'd29363};
                15'd4798 : data_rom <= {16'd14547, 16'd29361};
                15'd4799 : data_rom <= {16'd14550, 16'd29360};
                15'd4800 : data_rom <= {16'd14552, 16'd29359};
                15'd4801 : data_rom <= {16'd14555, 16'd29357};
                15'd4802 : data_rom <= {16'd14558, 16'd29356};
                15'd4803 : data_rom <= {16'd14561, 16'd29354};
                15'd4804 : data_rom <= {16'd14564, 16'd29353};
                15'd4805 : data_rom <= {16'd14567, 16'd29352};
                15'd4806 : data_rom <= {16'd14569, 16'd29350};
                15'd4807 : data_rom <= {16'd14572, 16'd29349};
                15'd4808 : data_rom <= {16'd14575, 16'd29347};
                15'd4809 : data_rom <= {16'd14578, 16'd29346};
                15'd4810 : data_rom <= {16'd14581, 16'd29345};
                15'd4811 : data_rom <= {16'd14583, 16'd29343};
                15'd4812 : data_rom <= {16'd14586, 16'd29342};
                15'd4813 : data_rom <= {16'd14589, 16'd29340};
                15'd4814 : data_rom <= {16'd14592, 16'd29339};
                15'd4815 : data_rom <= {16'd14595, 16'd29338};
                15'd4816 : data_rom <= {16'd14598, 16'd29336};
                15'd4817 : data_rom <= {16'd14600, 16'd29335};
                15'd4818 : data_rom <= {16'd14603, 16'd29333};
                15'd4819 : data_rom <= {16'd14606, 16'd29332};
                15'd4820 : data_rom <= {16'd14609, 16'd29331};
                15'd4821 : data_rom <= {16'd14612, 16'd29329};
                15'd4822 : data_rom <= {16'd14614, 16'd29328};
                15'd4823 : data_rom <= {16'd14617, 16'd29326};
                15'd4824 : data_rom <= {16'd14620, 16'd29325};
                15'd4825 : data_rom <= {16'd14623, 16'd29324};
                15'd4826 : data_rom <= {16'd14626, 16'd29322};
                15'd4827 : data_rom <= {16'd14628, 16'd29321};
                15'd4828 : data_rom <= {16'd14631, 16'd29319};
                15'd4829 : data_rom <= {16'd14634, 16'd29318};
                15'd4830 : data_rom <= {16'd14637, 16'd29317};
                15'd4831 : data_rom <= {16'd14640, 16'd29315};
                15'd4832 : data_rom <= {16'd14642, 16'd29314};
                15'd4833 : data_rom <= {16'd14645, 16'd29312};
                15'd4834 : data_rom <= {16'd14648, 16'd29311};
                15'd4835 : data_rom <= {16'd14651, 16'd29310};
                15'd4836 : data_rom <= {16'd14654, 16'd29308};
                15'd4837 : data_rom <= {16'd14657, 16'd29307};
                15'd4838 : data_rom <= {16'd14659, 16'd29305};
                15'd4839 : data_rom <= {16'd14662, 16'd29304};
                15'd4840 : data_rom <= {16'd14665, 16'd29303};
                15'd4841 : data_rom <= {16'd14668, 16'd29301};
                15'd4842 : data_rom <= {16'd14671, 16'd29300};
                15'd4843 : data_rom <= {16'd14673, 16'd29298};
                15'd4844 : data_rom <= {16'd14676, 16'd29297};
                15'd4845 : data_rom <= {16'd14679, 16'd29295};
                15'd4846 : data_rom <= {16'd14682, 16'd29294};
                15'd4847 : data_rom <= {16'd14685, 16'd29293};
                15'd4848 : data_rom <= {16'd14687, 16'd29291};
                15'd4849 : data_rom <= {16'd14690, 16'd29290};
                15'd4850 : data_rom <= {16'd14693, 16'd29288};
                15'd4851 : data_rom <= {16'd14696, 16'd29287};
                15'd4852 : data_rom <= {16'd14699, 16'd29286};
                15'd4853 : data_rom <= {16'd14701, 16'd29284};
                15'd4854 : data_rom <= {16'd14704, 16'd29283};
                15'd4855 : data_rom <= {16'd14707, 16'd29281};
                15'd4856 : data_rom <= {16'd14710, 16'd29280};
                15'd4857 : data_rom <= {16'd14713, 16'd29279};
                15'd4858 : data_rom <= {16'd14716, 16'd29277};
                15'd4859 : data_rom <= {16'd14718, 16'd29276};
                15'd4860 : data_rom <= {16'd14721, 16'd29274};
                15'd4861 : data_rom <= {16'd14724, 16'd29273};
                15'd4862 : data_rom <= {16'd14727, 16'd29272};
                15'd4863 : data_rom <= {16'd14730, 16'd29270};
                15'd4864 : data_rom <= {16'd14732, 16'd29269};
                15'd4865 : data_rom <= {16'd14735, 16'd29267};
                15'd4866 : data_rom <= {16'd14738, 16'd29266};
                15'd4867 : data_rom <= {16'd14741, 16'd29264};
                15'd4868 : data_rom <= {16'd14744, 16'd29263};
                15'd4869 : data_rom <= {16'd14746, 16'd29262};
                15'd4870 : data_rom <= {16'd14749, 16'd29260};
                15'd4871 : data_rom <= {16'd14752, 16'd29259};
                15'd4872 : data_rom <= {16'd14755, 16'd29257};
                15'd4873 : data_rom <= {16'd14758, 16'd29256};
                15'd4874 : data_rom <= {16'd14760, 16'd29255};
                15'd4875 : data_rom <= {16'd14763, 16'd29253};
                15'd4876 : data_rom <= {16'd14766, 16'd29252};
                15'd4877 : data_rom <= {16'd14769, 16'd29250};
                15'd4878 : data_rom <= {16'd14772, 16'd29249};
                15'd4879 : data_rom <= {16'd14774, 16'd29247};
                15'd4880 : data_rom <= {16'd14777, 16'd29246};
                15'd4881 : data_rom <= {16'd14780, 16'd29245};
                15'd4882 : data_rom <= {16'd14783, 16'd29243};
                15'd4883 : data_rom <= {16'd14786, 16'd29242};
                15'd4884 : data_rom <= {16'd14788, 16'd29240};
                15'd4885 : data_rom <= {16'd14791, 16'd29239};
                15'd4886 : data_rom <= {16'd14794, 16'd29238};
                15'd4887 : data_rom <= {16'd14797, 16'd29236};
                15'd4888 : data_rom <= {16'd14800, 16'd29235};
                15'd4889 : data_rom <= {16'd14802, 16'd29233};
                15'd4890 : data_rom <= {16'd14805, 16'd29232};
                15'd4891 : data_rom <= {16'd14808, 16'd29230};
                15'd4892 : data_rom <= {16'd14811, 16'd29229};
                15'd4893 : data_rom <= {16'd14814, 16'd29228};
                15'd4894 : data_rom <= {16'd14816, 16'd29226};
                15'd4895 : data_rom <= {16'd14819, 16'd29225};
                15'd4896 : data_rom <= {16'd14822, 16'd29223};
                15'd4897 : data_rom <= {16'd14825, 16'd29222};
                15'd4898 : data_rom <= {16'd14828, 16'd29221};
                15'd4899 : data_rom <= {16'd14830, 16'd29219};
                15'd4900 : data_rom <= {16'd14833, 16'd29218};
                15'd4901 : data_rom <= {16'd14836, 16'd29216};
                15'd4902 : data_rom <= {16'd14839, 16'd29215};
                15'd4903 : data_rom <= {16'd14842, 16'd29213};
                15'd4904 : data_rom <= {16'd14844, 16'd29212};
                15'd4905 : data_rom <= {16'd14847, 16'd29211};
                15'd4906 : data_rom <= {16'd14850, 16'd29209};
                15'd4907 : data_rom <= {16'd14853, 16'd29208};
                15'd4908 : data_rom <= {16'd14856, 16'd29206};
                15'd4909 : data_rom <= {16'd14858, 16'd29205};
                15'd4910 : data_rom <= {16'd14861, 16'd29203};
                15'd4911 : data_rom <= {16'd14864, 16'd29202};
                15'd4912 : data_rom <= {16'd14867, 16'd29201};
                15'd4913 : data_rom <= {16'd14870, 16'd29199};
                15'd4914 : data_rom <= {16'd14872, 16'd29198};
                15'd4915 : data_rom <= {16'd14875, 16'd29196};
                15'd4916 : data_rom <= {16'd14878, 16'd29195};
                15'd4917 : data_rom <= {16'd14881, 16'd29193};
                15'd4918 : data_rom <= {16'd14884, 16'd29192};
                15'd4919 : data_rom <= {16'd14886, 16'd29191};
                15'd4920 : data_rom <= {16'd14889, 16'd29189};
                15'd4921 : data_rom <= {16'd14892, 16'd29188};
                15'd4922 : data_rom <= {16'd14895, 16'd29186};
                15'd4923 : data_rom <= {16'd14898, 16'd29185};
                15'd4924 : data_rom <= {16'd14900, 16'd29183};
                15'd4925 : data_rom <= {16'd14903, 16'd29182};
                15'd4926 : data_rom <= {16'd14906, 16'd29181};
                15'd4927 : data_rom <= {16'd14909, 16'd29179};
                15'd4928 : data_rom <= {16'd14912, 16'd29178};
                15'd4929 : data_rom <= {16'd14914, 16'd29176};
                15'd4930 : data_rom <= {16'd14917, 16'd29175};
                15'd4931 : data_rom <= {16'd14920, 16'd29173};
                15'd4932 : data_rom <= {16'd14923, 16'd29172};
                15'd4933 : data_rom <= {16'd14926, 16'd29171};
                15'd4934 : data_rom <= {16'd14928, 16'd29169};
                15'd4935 : data_rom <= {16'd14931, 16'd29168};
                15'd4936 : data_rom <= {16'd14934, 16'd29166};
                15'd4937 : data_rom <= {16'd14937, 16'd29165};
                15'd4938 : data_rom <= {16'd14940, 16'd29163};
                15'd4939 : data_rom <= {16'd14942, 16'd29162};
                15'd4940 : data_rom <= {16'd14945, 16'd29161};
                15'd4941 : data_rom <= {16'd14948, 16'd29159};
                15'd4942 : data_rom <= {16'd14951, 16'd29158};
                15'd4943 : data_rom <= {16'd14954, 16'd29156};
                15'd4944 : data_rom <= {16'd14956, 16'd29155};
                15'd4945 : data_rom <= {16'd14959, 16'd29153};
                15'd4946 : data_rom <= {16'd14962, 16'd29152};
                15'd4947 : data_rom <= {16'd14965, 16'd29151};
                15'd4948 : data_rom <= {16'd14968, 16'd29149};
                15'd4949 : data_rom <= {16'd14970, 16'd29148};
                15'd4950 : data_rom <= {16'd14973, 16'd29146};
                15'd4951 : data_rom <= {16'd14976, 16'd29145};
                15'd4952 : data_rom <= {16'd14979, 16'd29143};
                15'd4953 : data_rom <= {16'd14982, 16'd29142};
                15'd4954 : data_rom <= {16'd14984, 16'd29140};
                15'd4955 : data_rom <= {16'd14987, 16'd29139};
                15'd4956 : data_rom <= {16'd14990, 16'd29138};
                15'd4957 : data_rom <= {16'd14993, 16'd29136};
                15'd4958 : data_rom <= {16'd14996, 16'd29135};
                15'd4959 : data_rom <= {16'd14998, 16'd29133};
                15'd4960 : data_rom <= {16'd15001, 16'd29132};
                15'd4961 : data_rom <= {16'd15004, 16'd29130};
                15'd4962 : data_rom <= {16'd15007, 16'd29129};
                15'd4963 : data_rom <= {16'd15009, 16'd29128};
                15'd4964 : data_rom <= {16'd15012, 16'd29126};
                15'd4965 : data_rom <= {16'd15015, 16'd29125};
                15'd4966 : data_rom <= {16'd15018, 16'd29123};
                15'd4967 : data_rom <= {16'd15021, 16'd29122};
                15'd4968 : data_rom <= {16'd15023, 16'd29120};
                15'd4969 : data_rom <= {16'd15026, 16'd29119};
                15'd4970 : data_rom <= {16'd15029, 16'd29117};
                15'd4971 : data_rom <= {16'd15032, 16'd29116};
                15'd4972 : data_rom <= {16'd15035, 16'd29115};
                15'd4973 : data_rom <= {16'd15037, 16'd29113};
                15'd4974 : data_rom <= {16'd15040, 16'd29112};
                15'd4975 : data_rom <= {16'd15043, 16'd29110};
                15'd4976 : data_rom <= {16'd15046, 16'd29109};
                15'd4977 : data_rom <= {16'd15049, 16'd29107};
                15'd4978 : data_rom <= {16'd15051, 16'd29106};
                15'd4979 : data_rom <= {16'd15054, 16'd29104};
                15'd4980 : data_rom <= {16'd15057, 16'd29103};
                15'd4981 : data_rom <= {16'd15060, 16'd29102};
                15'd4982 : data_rom <= {16'd15063, 16'd29100};
                15'd4983 : data_rom <= {16'd15065, 16'd29099};
                15'd4984 : data_rom <= {16'd15068, 16'd29097};
                15'd4985 : data_rom <= {16'd15071, 16'd29096};
                15'd4986 : data_rom <= {16'd15074, 16'd29094};
                15'd4987 : data_rom <= {16'd15076, 16'd29093};
                15'd4988 : data_rom <= {16'd15079, 16'd29091};
                15'd4989 : data_rom <= {16'd15082, 16'd29090};
                15'd4990 : data_rom <= {16'd15085, 16'd29089};
                15'd4991 : data_rom <= {16'd15088, 16'd29087};
                15'd4992 : data_rom <= {16'd15090, 16'd29086};
                15'd4993 : data_rom <= {16'd15093, 16'd29084};
                15'd4994 : data_rom <= {16'd15096, 16'd29083};
                15'd4995 : data_rom <= {16'd15099, 16'd29081};
                15'd4996 : data_rom <= {16'd15102, 16'd29080};
                15'd4997 : data_rom <= {16'd15104, 16'd29078};
                15'd4998 : data_rom <= {16'd15107, 16'd29077};
                15'd4999 : data_rom <= {16'd15110, 16'd29076};
                15'd5000 : data_rom <= {16'd15113, 16'd29074};
                15'd5001 : data_rom <= {16'd15116, 16'd29073};
                15'd5002 : data_rom <= {16'd15118, 16'd29071};
                15'd5003 : data_rom <= {16'd15121, 16'd29070};
                15'd5004 : data_rom <= {16'd15124, 16'd29068};
                15'd5005 : data_rom <= {16'd15127, 16'd29067};
                15'd5006 : data_rom <= {16'd15129, 16'd29065};
                15'd5007 : data_rom <= {16'd15132, 16'd29064};
                15'd5008 : data_rom <= {16'd15135, 16'd29062};
                15'd5009 : data_rom <= {16'd15138, 16'd29061};
                15'd5010 : data_rom <= {16'd15141, 16'd29060};
                15'd5011 : data_rom <= {16'd15143, 16'd29058};
                15'd5012 : data_rom <= {16'd15146, 16'd29057};
                15'd5013 : data_rom <= {16'd15149, 16'd29055};
                15'd5014 : data_rom <= {16'd15152, 16'd29054};
                15'd5015 : data_rom <= {16'd15155, 16'd29052};
                15'd5016 : data_rom <= {16'd15157, 16'd29051};
                15'd5017 : data_rom <= {16'd15160, 16'd29049};
                15'd5018 : data_rom <= {16'd15163, 16'd29048};
                15'd5019 : data_rom <= {16'd15166, 16'd29047};
                15'd5020 : data_rom <= {16'd15168, 16'd29045};
                15'd5021 : data_rom <= {16'd15171, 16'd29044};
                15'd5022 : data_rom <= {16'd15174, 16'd29042};
                15'd5023 : data_rom <= {16'd15177, 16'd29041};
                15'd5024 : data_rom <= {16'd15180, 16'd29039};
                15'd5025 : data_rom <= {16'd15182, 16'd29038};
                15'd5026 : data_rom <= {16'd15185, 16'd29036};
                15'd5027 : data_rom <= {16'd15188, 16'd29035};
                15'd5028 : data_rom <= {16'd15191, 16'd29033};
                15'd5029 : data_rom <= {16'd15194, 16'd29032};
                15'd5030 : data_rom <= {16'd15196, 16'd29031};
                15'd5031 : data_rom <= {16'd15199, 16'd29029};
                15'd5032 : data_rom <= {16'd15202, 16'd29028};
                15'd5033 : data_rom <= {16'd15205, 16'd29026};
                15'd5034 : data_rom <= {16'd15207, 16'd29025};
                15'd5035 : data_rom <= {16'd15210, 16'd29023};
                15'd5036 : data_rom <= {16'd15213, 16'd29022};
                15'd5037 : data_rom <= {16'd15216, 16'd29020};
                15'd5038 : data_rom <= {16'd15219, 16'd29019};
                15'd5039 : data_rom <= {16'd15221, 16'd29017};
                15'd5040 : data_rom <= {16'd15224, 16'd29016};
                15'd5041 : data_rom <= {16'd15227, 16'd29014};
                15'd5042 : data_rom <= {16'd15230, 16'd29013};
                15'd5043 : data_rom <= {16'd15232, 16'd29012};
                15'd5044 : data_rom <= {16'd15235, 16'd29010};
                15'd5045 : data_rom <= {16'd15238, 16'd29009};
                15'd5046 : data_rom <= {16'd15241, 16'd29007};
                15'd5047 : data_rom <= {16'd15244, 16'd29006};
                15'd5048 : data_rom <= {16'd15246, 16'd29004};
                15'd5049 : data_rom <= {16'd15249, 16'd29003};
                15'd5050 : data_rom <= {16'd15252, 16'd29001};
                15'd5051 : data_rom <= {16'd15255, 16'd29000};
                15'd5052 : data_rom <= {16'd15257, 16'd28998};
                15'd5053 : data_rom <= {16'd15260, 16'd28997};
                15'd5054 : data_rom <= {16'd15263, 16'd28995};
                15'd5055 : data_rom <= {16'd15266, 16'd28994};
                15'd5056 : data_rom <= {16'd15269, 16'd28993};
                15'd5057 : data_rom <= {16'd15271, 16'd28991};
                15'd5058 : data_rom <= {16'd15274, 16'd28990};
                15'd5059 : data_rom <= {16'd15277, 16'd28988};
                15'd5060 : data_rom <= {16'd15280, 16'd28987};
                15'd5061 : data_rom <= {16'd15283, 16'd28985};
                15'd5062 : data_rom <= {16'd15285, 16'd28984};
                15'd5063 : data_rom <= {16'd15288, 16'd28982};
                15'd5064 : data_rom <= {16'd15291, 16'd28981};
                15'd5065 : data_rom <= {16'd15294, 16'd28979};
                15'd5066 : data_rom <= {16'd15296, 16'd28978};
                15'd5067 : data_rom <= {16'd15299, 16'd28976};
                15'd5068 : data_rom <= {16'd15302, 16'd28975};
                15'd5069 : data_rom <= {16'd15305, 16'd28973};
                15'd5070 : data_rom <= {16'd15308, 16'd28972};
                15'd5071 : data_rom <= {16'd15310, 16'd28971};
                15'd5072 : data_rom <= {16'd15313, 16'd28969};
                15'd5073 : data_rom <= {16'd15316, 16'd28968};
                15'd5074 : data_rom <= {16'd15319, 16'd28966};
                15'd5075 : data_rom <= {16'd15321, 16'd28965};
                15'd5076 : data_rom <= {16'd15324, 16'd28963};
                15'd5077 : data_rom <= {16'd15327, 16'd28962};
                15'd5078 : data_rom <= {16'd15330, 16'd28960};
                15'd5079 : data_rom <= {16'd15332, 16'd28959};
                15'd5080 : data_rom <= {16'd15335, 16'd28957};
                15'd5081 : data_rom <= {16'd15338, 16'd28956};
                15'd5082 : data_rom <= {16'd15341, 16'd28954};
                15'd5083 : data_rom <= {16'd15344, 16'd28953};
                15'd5084 : data_rom <= {16'd15346, 16'd28951};
                15'd5085 : data_rom <= {16'd15349, 16'd28950};
                15'd5086 : data_rom <= {16'd15352, 16'd28949};
                15'd5087 : data_rom <= {16'd15355, 16'd28947};
                15'd5088 : data_rom <= {16'd15357, 16'd28946};
                15'd5089 : data_rom <= {16'd15360, 16'd28944};
                15'd5090 : data_rom <= {16'd15363, 16'd28943};
                15'd5091 : data_rom <= {16'd15366, 16'd28941};
                15'd5092 : data_rom <= {16'd15369, 16'd28940};
                15'd5093 : data_rom <= {16'd15371, 16'd28938};
                15'd5094 : data_rom <= {16'd15374, 16'd28937};
                15'd5095 : data_rom <= {16'd15377, 16'd28935};
                15'd5096 : data_rom <= {16'd15380, 16'd28934};
                15'd5097 : data_rom <= {16'd15382, 16'd28932};
                15'd5098 : data_rom <= {16'd15385, 16'd28931};
                15'd5099 : data_rom <= {16'd15388, 16'd28929};
                15'd5100 : data_rom <= {16'd15391, 16'd28928};
                15'd5101 : data_rom <= {16'd15394, 16'd28926};
                15'd5102 : data_rom <= {16'd15396, 16'd28925};
                15'd5103 : data_rom <= {16'd15399, 16'd28923};
                15'd5104 : data_rom <= {16'd15402, 16'd28922};
                15'd5105 : data_rom <= {16'd15405, 16'd28920};
                15'd5106 : data_rom <= {16'd15407, 16'd28919};
                15'd5107 : data_rom <= {16'd15410, 16'd28918};
                15'd5108 : data_rom <= {16'd15413, 16'd28916};
                15'd5109 : data_rom <= {16'd15416, 16'd28915};
                15'd5110 : data_rom <= {16'd15419, 16'd28913};
                15'd5111 : data_rom <= {16'd15421, 16'd28912};
                15'd5112 : data_rom <= {16'd15424, 16'd28910};
                15'd5113 : data_rom <= {16'd15427, 16'd28909};
                15'd5114 : data_rom <= {16'd15430, 16'd28907};
                15'd5115 : data_rom <= {16'd15432, 16'd28906};
                15'd5116 : data_rom <= {16'd15435, 16'd28904};
                15'd5117 : data_rom <= {16'd15438, 16'd28903};
                15'd5118 : data_rom <= {16'd15441, 16'd28901};
                15'd5119 : data_rom <= {16'd15443, 16'd28900};
                15'd5120 : data_rom <= {16'd15446, 16'd28898};
                15'd5121 : data_rom <= {16'd15449, 16'd28897};
                15'd5122 : data_rom <= {16'd15452, 16'd28895};
                15'd5123 : data_rom <= {16'd15455, 16'd28894};
                15'd5124 : data_rom <= {16'd15457, 16'd28892};
                15'd5125 : data_rom <= {16'd15460, 16'd28891};
                15'd5126 : data_rom <= {16'd15463, 16'd28889};
                15'd5127 : data_rom <= {16'd15466, 16'd28888};
                15'd5128 : data_rom <= {16'd15468, 16'd28886};
                15'd5129 : data_rom <= {16'd15471, 16'd28885};
                15'd5130 : data_rom <= {16'd15474, 16'd28883};
                15'd5131 : data_rom <= {16'd15477, 16'd28882};
                15'd5132 : data_rom <= {16'd15479, 16'd28881};
                15'd5133 : data_rom <= {16'd15482, 16'd28879};
                15'd5134 : data_rom <= {16'd15485, 16'd28878};
                15'd5135 : data_rom <= {16'd15488, 16'd28876};
                15'd5136 : data_rom <= {16'd15491, 16'd28875};
                15'd5137 : data_rom <= {16'd15493, 16'd28873};
                15'd5138 : data_rom <= {16'd15496, 16'd28872};
                15'd5139 : data_rom <= {16'd15499, 16'd28870};
                15'd5140 : data_rom <= {16'd15502, 16'd28869};
                15'd5141 : data_rom <= {16'd15504, 16'd28867};
                15'd5142 : data_rom <= {16'd15507, 16'd28866};
                15'd5143 : data_rom <= {16'd15510, 16'd28864};
                15'd5144 : data_rom <= {16'd15513, 16'd28863};
                15'd5145 : data_rom <= {16'd15515, 16'd28861};
                15'd5146 : data_rom <= {16'd15518, 16'd28860};
                15'd5147 : data_rom <= {16'd15521, 16'd28858};
                15'd5148 : data_rom <= {16'd15524, 16'd28857};
                15'd5149 : data_rom <= {16'd15527, 16'd28855};
                15'd5150 : data_rom <= {16'd15529, 16'd28854};
                15'd5151 : data_rom <= {16'd15532, 16'd28852};
                15'd5152 : data_rom <= {16'd15535, 16'd28851};
                15'd5153 : data_rom <= {16'd15538, 16'd28849};
                15'd5154 : data_rom <= {16'd15540, 16'd28848};
                15'd5155 : data_rom <= {16'd15543, 16'd28846};
                15'd5156 : data_rom <= {16'd15546, 16'd28845};
                15'd5157 : data_rom <= {16'd15549, 16'd28843};
                15'd5158 : data_rom <= {16'd15551, 16'd28842};
                15'd5159 : data_rom <= {16'd15554, 16'd28840};
                15'd5160 : data_rom <= {16'd15557, 16'd28839};
                15'd5161 : data_rom <= {16'd15560, 16'd28837};
                15'd5162 : data_rom <= {16'd15562, 16'd28836};
                15'd5163 : data_rom <= {16'd15565, 16'd28834};
                15'd5164 : data_rom <= {16'd15568, 16'd28833};
                15'd5165 : data_rom <= {16'd15571, 16'd28831};
                15'd5166 : data_rom <= {16'd15574, 16'd28830};
                15'd5167 : data_rom <= {16'd15576, 16'd28828};
                15'd5168 : data_rom <= {16'd15579, 16'd28827};
                15'd5169 : data_rom <= {16'd15582, 16'd28825};
                15'd5170 : data_rom <= {16'd15585, 16'd28824};
                15'd5171 : data_rom <= {16'd15587, 16'd28822};
                15'd5172 : data_rom <= {16'd15590, 16'd28821};
                15'd5173 : data_rom <= {16'd15593, 16'd28819};
                15'd5174 : data_rom <= {16'd15596, 16'd28818};
                15'd5175 : data_rom <= {16'd15598, 16'd28816};
                15'd5176 : data_rom <= {16'd15601, 16'd28815};
                15'd5177 : data_rom <= {16'd15604, 16'd28813};
                15'd5178 : data_rom <= {16'd15607, 16'd28812};
                15'd5179 : data_rom <= {16'd15609, 16'd28810};
                15'd5180 : data_rom <= {16'd15612, 16'd28809};
                15'd5181 : data_rom <= {16'd15615, 16'd28807};
                15'd5182 : data_rom <= {16'd15618, 16'd28806};
                15'd5183 : data_rom <= {16'd15620, 16'd28804};
                15'd5184 : data_rom <= {16'd15623, 16'd28803};
                15'd5185 : data_rom <= {16'd15626, 16'd28801};
                15'd5186 : data_rom <= {16'd15629, 16'd28800};
                15'd5187 : data_rom <= {16'd15632, 16'd28798};
                15'd5188 : data_rom <= {16'd15634, 16'd28797};
                15'd5189 : data_rom <= {16'd15637, 16'd28795};
                15'd5190 : data_rom <= {16'd15640, 16'd28794};
                15'd5191 : data_rom <= {16'd15643, 16'd28792};
                15'd5192 : data_rom <= {16'd15645, 16'd28791};
                15'd5193 : data_rom <= {16'd15648, 16'd28789};
                15'd5194 : data_rom <= {16'd15651, 16'd28788};
                15'd5195 : data_rom <= {16'd15654, 16'd28786};
                15'd5196 : data_rom <= {16'd15656, 16'd28785};
                15'd5197 : data_rom <= {16'd15659, 16'd28783};
                15'd5198 : data_rom <= {16'd15662, 16'd28782};
                15'd5199 : data_rom <= {16'd15665, 16'd28780};
                15'd5200 : data_rom <= {16'd15667, 16'd28779};
                15'd5201 : data_rom <= {16'd15670, 16'd28777};
                15'd5202 : data_rom <= {16'd15673, 16'd28776};
                15'd5203 : data_rom <= {16'd15676, 16'd28774};
                15'd5204 : data_rom <= {16'd15678, 16'd28773};
                15'd5205 : data_rom <= {16'd15681, 16'd28771};
                15'd5206 : data_rom <= {16'd15684, 16'd28770};
                15'd5207 : data_rom <= {16'd15687, 16'd28768};
                15'd5208 : data_rom <= {16'd15689, 16'd28767};
                15'd5209 : data_rom <= {16'd15692, 16'd28765};
                15'd5210 : data_rom <= {16'd15695, 16'd28764};
                15'd5211 : data_rom <= {16'd15698, 16'd28762};
                15'd5212 : data_rom <= {16'd15701, 16'd28761};
                15'd5213 : data_rom <= {16'd15703, 16'd28759};
                15'd5214 : data_rom <= {16'd15706, 16'd28758};
                15'd5215 : data_rom <= {16'd15709, 16'd28756};
                15'd5216 : data_rom <= {16'd15712, 16'd28755};
                15'd5217 : data_rom <= {16'd15714, 16'd28753};
                15'd5218 : data_rom <= {16'd15717, 16'd28752};
                15'd5219 : data_rom <= {16'd15720, 16'd28750};
                15'd5220 : data_rom <= {16'd15723, 16'd28749};
                15'd5221 : data_rom <= {16'd15725, 16'd28747};
                15'd5222 : data_rom <= {16'd15728, 16'd28746};
                15'd5223 : data_rom <= {16'd15731, 16'd28744};
                15'd5224 : data_rom <= {16'd15734, 16'd28743};
                15'd5225 : data_rom <= {16'd15736, 16'd28741};
                15'd5226 : data_rom <= {16'd15739, 16'd28740};
                15'd5227 : data_rom <= {16'd15742, 16'd28738};
                15'd5228 : data_rom <= {16'd15745, 16'd28737};
                15'd5229 : data_rom <= {16'd15747, 16'd28735};
                15'd5230 : data_rom <= {16'd15750, 16'd28734};
                15'd5231 : data_rom <= {16'd15753, 16'd28732};
                15'd5232 : data_rom <= {16'd15756, 16'd28731};
                15'd5233 : data_rom <= {16'd15758, 16'd28729};
                15'd5234 : data_rom <= {16'd15761, 16'd28728};
                15'd5235 : data_rom <= {16'd15764, 16'd28726};
                15'd5236 : data_rom <= {16'd15767, 16'd28725};
                15'd5237 : data_rom <= {16'd15769, 16'd28723};
                15'd5238 : data_rom <= {16'd15772, 16'd28722};
                15'd5239 : data_rom <= {16'd15775, 16'd28720};
                15'd5240 : data_rom <= {16'd15778, 16'd28719};
                15'd5241 : data_rom <= {16'd15780, 16'd28717};
                15'd5242 : data_rom <= {16'd15783, 16'd28716};
                15'd5243 : data_rom <= {16'd15786, 16'd28714};
                15'd5244 : data_rom <= {16'd15789, 16'd28713};
                15'd5245 : data_rom <= {16'd15791, 16'd28711};
                15'd5246 : data_rom <= {16'd15794, 16'd28710};
                15'd5247 : data_rom <= {16'd15797, 16'd28708};
                15'd5248 : data_rom <= {16'd15800, 16'd28707};
                15'd5249 : data_rom <= {16'd15802, 16'd28705};
                15'd5250 : data_rom <= {16'd15805, 16'd28704};
                15'd5251 : data_rom <= {16'd15808, 16'd28702};
                15'd5252 : data_rom <= {16'd15811, 16'd28701};
                15'd5253 : data_rom <= {16'd15813, 16'd28699};
                15'd5254 : data_rom <= {16'd15816, 16'd28697};
                15'd5255 : data_rom <= {16'd15819, 16'd28696};
                15'd5256 : data_rom <= {16'd15822, 16'd28694};
                15'd5257 : data_rom <= {16'd15824, 16'd28693};
                15'd5258 : data_rom <= {16'd15827, 16'd28691};
                15'd5259 : data_rom <= {16'd15830, 16'd28690};
                15'd5260 : data_rom <= {16'd15833, 16'd28688};
                15'd5261 : data_rom <= {16'd15835, 16'd28687};
                15'd5262 : data_rom <= {16'd15838, 16'd28685};
                15'd5263 : data_rom <= {16'd15841, 16'd28684};
                15'd5264 : data_rom <= {16'd15844, 16'd28682};
                15'd5265 : data_rom <= {16'd15846, 16'd28681};
                15'd5266 : data_rom <= {16'd15849, 16'd28679};
                15'd5267 : data_rom <= {16'd15852, 16'd28678};
                15'd5268 : data_rom <= {16'd15855, 16'd28676};
                15'd5269 : data_rom <= {16'd15857, 16'd28675};
                15'd5270 : data_rom <= {16'd15860, 16'd28673};
                15'd5271 : data_rom <= {16'd15863, 16'd28672};
                15'd5272 : data_rom <= {16'd15866, 16'd28670};
                15'd5273 : data_rom <= {16'd15868, 16'd28669};
                15'd5274 : data_rom <= {16'd15871, 16'd28667};
                15'd5275 : data_rom <= {16'd15874, 16'd28666};
                15'd5276 : data_rom <= {16'd15877, 16'd28664};
                15'd5277 : data_rom <= {16'd15879, 16'd28663};
                15'd5278 : data_rom <= {16'd15882, 16'd28661};
                15'd5279 : data_rom <= {16'd15885, 16'd28659};
                15'd5280 : data_rom <= {16'd15888, 16'd28658};
                15'd5281 : data_rom <= {16'd15890, 16'd28656};
                15'd5282 : data_rom <= {16'd15893, 16'd28655};
                15'd5283 : data_rom <= {16'd15896, 16'd28653};
                15'd5284 : data_rom <= {16'd15899, 16'd28652};
                15'd5285 : data_rom <= {16'd15901, 16'd28650};
                15'd5286 : data_rom <= {16'd15904, 16'd28649};
                15'd5287 : data_rom <= {16'd15907, 16'd28647};
                15'd5288 : data_rom <= {16'd15910, 16'd28646};
                15'd5289 : data_rom <= {16'd15912, 16'd28644};
                15'd5290 : data_rom <= {16'd15915, 16'd28643};
                15'd5291 : data_rom <= {16'd15918, 16'd28641};
                15'd5292 : data_rom <= {16'd15921, 16'd28640};
                15'd5293 : data_rom <= {16'd15923, 16'd28638};
                15'd5294 : data_rom <= {16'd15926, 16'd28637};
                15'd5295 : data_rom <= {16'd15929, 16'd28635};
                15'd5296 : data_rom <= {16'd15932, 16'd28634};
                15'd5297 : data_rom <= {16'd15934, 16'd28632};
                15'd5298 : data_rom <= {16'd15937, 16'd28631};
                15'd5299 : data_rom <= {16'd15940, 16'd28629};
                15'd5300 : data_rom <= {16'd15943, 16'd28627};
                15'd5301 : data_rom <= {16'd15945, 16'd28626};
                15'd5302 : data_rom <= {16'd15948, 16'd28624};
                15'd5303 : data_rom <= {16'd15951, 16'd28623};
                15'd5304 : data_rom <= {16'd15954, 16'd28621};
                15'd5305 : data_rom <= {16'd15956, 16'd28620};
                15'd5306 : data_rom <= {16'd15959, 16'd28618};
                15'd5307 : data_rom <= {16'd15962, 16'd28617};
                15'd5308 : data_rom <= {16'd15965, 16'd28615};
                15'd5309 : data_rom <= {16'd15967, 16'd28614};
                15'd5310 : data_rom <= {16'd15970, 16'd28612};
                15'd5311 : data_rom <= {16'd15973, 16'd28611};
                15'd5312 : data_rom <= {16'd15976, 16'd28609};
                15'd5313 : data_rom <= {16'd15978, 16'd28608};
                15'd5314 : data_rom <= {16'd15981, 16'd28606};
                15'd5315 : data_rom <= {16'd15984, 16'd28604};
                15'd5316 : data_rom <= {16'd15987, 16'd28603};
                15'd5317 : data_rom <= {16'd15989, 16'd28601};
                15'd5318 : data_rom <= {16'd15992, 16'd28600};
                15'd5319 : data_rom <= {16'd15995, 16'd28598};
                15'd5320 : data_rom <= {16'd15997, 16'd28597};
                15'd5321 : data_rom <= {16'd16000, 16'd28595};
                15'd5322 : data_rom <= {16'd16003, 16'd28594};
                15'd5323 : data_rom <= {16'd16006, 16'd28592};
                15'd5324 : data_rom <= {16'd16008, 16'd28591};
                15'd5325 : data_rom <= {16'd16011, 16'd28589};
                15'd5326 : data_rom <= {16'd16014, 16'd28588};
                15'd5327 : data_rom <= {16'd16017, 16'd28586};
                15'd5328 : data_rom <= {16'd16019, 16'd28585};
                15'd5329 : data_rom <= {16'd16022, 16'd28583};
                15'd5330 : data_rom <= {16'd16025, 16'd28581};
                15'd5331 : data_rom <= {16'd16028, 16'd28580};
                15'd5332 : data_rom <= {16'd16030, 16'd28578};
                15'd5333 : data_rom <= {16'd16033, 16'd28577};
                15'd5334 : data_rom <= {16'd16036, 16'd28575};
                15'd5335 : data_rom <= {16'd16039, 16'd28574};
                15'd5336 : data_rom <= {16'd16041, 16'd28572};
                15'd5337 : data_rom <= {16'd16044, 16'd28571};
                15'd5338 : data_rom <= {16'd16047, 16'd28569};
                15'd5339 : data_rom <= {16'd16050, 16'd28568};
                15'd5340 : data_rom <= {16'd16052, 16'd28566};
                15'd5341 : data_rom <= {16'd16055, 16'd28565};
                15'd5342 : data_rom <= {16'd16058, 16'd28563};
                15'd5343 : data_rom <= {16'd16060, 16'd28561};
                15'd5344 : data_rom <= {16'd16063, 16'd28560};
                15'd5345 : data_rom <= {16'd16066, 16'd28558};
                15'd5346 : data_rom <= {16'd16069, 16'd28557};
                15'd5347 : data_rom <= {16'd16071, 16'd28555};
                15'd5348 : data_rom <= {16'd16074, 16'd28554};
                15'd5349 : data_rom <= {16'd16077, 16'd28552};
                15'd5350 : data_rom <= {16'd16080, 16'd28551};
                15'd5351 : data_rom <= {16'd16082, 16'd28549};
                15'd5352 : data_rom <= {16'd16085, 16'd28548};
                15'd5353 : data_rom <= {16'd16088, 16'd28546};
                15'd5354 : data_rom <= {16'd16091, 16'd28545};
                15'd5355 : data_rom <= {16'd16093, 16'd28543};
                15'd5356 : data_rom <= {16'd16096, 16'd28541};
                15'd5357 : data_rom <= {16'd16099, 16'd28540};
                15'd5358 : data_rom <= {16'd16102, 16'd28538};
                15'd5359 : data_rom <= {16'd16104, 16'd28537};
                15'd5360 : data_rom <= {16'd16107, 16'd28535};
                15'd5361 : data_rom <= {16'd16110, 16'd28534};
                15'd5362 : data_rom <= {16'd16112, 16'd28532};
                15'd5363 : data_rom <= {16'd16115, 16'd28531};
                15'd5364 : data_rom <= {16'd16118, 16'd28529};
                15'd5365 : data_rom <= {16'd16121, 16'd28528};
                15'd5366 : data_rom <= {16'd16123, 16'd28526};
                15'd5367 : data_rom <= {16'd16126, 16'd28524};
                15'd5368 : data_rom <= {16'd16129, 16'd28523};
                15'd5369 : data_rom <= {16'd16132, 16'd28521};
                15'd5370 : data_rom <= {16'd16134, 16'd28520};
                15'd5371 : data_rom <= {16'd16137, 16'd28518};
                15'd5372 : data_rom <= {16'd16140, 16'd28517};
                15'd5373 : data_rom <= {16'd16143, 16'd28515};
                15'd5374 : data_rom <= {16'd16145, 16'd28514};
                15'd5375 : data_rom <= {16'd16148, 16'd28512};
                15'd5376 : data_rom <= {16'd16151, 16'd28511};
                15'd5377 : data_rom <= {16'd16154, 16'd28509};
                15'd5378 : data_rom <= {16'd16156, 16'd28507};
                15'd5379 : data_rom <= {16'd16159, 16'd28506};
                15'd5380 : data_rom <= {16'd16162, 16'd28504};
                15'd5381 : data_rom <= {16'd16164, 16'd28503};
                15'd5382 : data_rom <= {16'd16167, 16'd28501};
                15'd5383 : data_rom <= {16'd16170, 16'd28500};
                15'd5384 : data_rom <= {16'd16173, 16'd28498};
                15'd5385 : data_rom <= {16'd16175, 16'd28497};
                15'd5386 : data_rom <= {16'd16178, 16'd28495};
                15'd5387 : data_rom <= {16'd16181, 16'd28493};
                15'd5388 : data_rom <= {16'd16184, 16'd28492};
                15'd5389 : data_rom <= {16'd16186, 16'd28490};
                15'd5390 : data_rom <= {16'd16189, 16'd28489};
                15'd5391 : data_rom <= {16'd16192, 16'd28487};
                15'd5392 : data_rom <= {16'd16194, 16'd28486};
                15'd5393 : data_rom <= {16'd16197, 16'd28484};
                15'd5394 : data_rom <= {16'd16200, 16'd28483};
                15'd5395 : data_rom <= {16'd16203, 16'd28481};
                15'd5396 : data_rom <= {16'd16205, 16'd28479};
                15'd5397 : data_rom <= {16'd16208, 16'd28478};
                15'd5398 : data_rom <= {16'd16211, 16'd28476};
                15'd5399 : data_rom <= {16'd16214, 16'd28475};
                15'd5400 : data_rom <= {16'd16216, 16'd28473};
                15'd5401 : data_rom <= {16'd16219, 16'd28472};
                15'd5402 : data_rom <= {16'd16222, 16'd28470};
                15'd5403 : data_rom <= {16'd16225, 16'd28469};
                15'd5404 : data_rom <= {16'd16227, 16'd28467};
                15'd5405 : data_rom <= {16'd16230, 16'd28466};
                15'd5406 : data_rom <= {16'd16233, 16'd28464};
                15'd5407 : data_rom <= {16'd16235, 16'd28462};
                15'd5408 : data_rom <= {16'd16238, 16'd28461};
                15'd5409 : data_rom <= {16'd16241, 16'd28459};
                15'd5410 : data_rom <= {16'd16244, 16'd28458};
                15'd5411 : data_rom <= {16'd16246, 16'd28456};
                15'd5412 : data_rom <= {16'd16249, 16'd28455};
                15'd5413 : data_rom <= {16'd16252, 16'd28453};
                15'd5414 : data_rom <= {16'd16255, 16'd28451};
                15'd5415 : data_rom <= {16'd16257, 16'd28450};
                15'd5416 : data_rom <= {16'd16260, 16'd28448};
                15'd5417 : data_rom <= {16'd16263, 16'd28447};
                15'd5418 : data_rom <= {16'd16265, 16'd28445};
                15'd5419 : data_rom <= {16'd16268, 16'd28444};
                15'd5420 : data_rom <= {16'd16271, 16'd28442};
                15'd5421 : data_rom <= {16'd16274, 16'd28441};
                15'd5422 : data_rom <= {16'd16276, 16'd28439};
                15'd5423 : data_rom <= {16'd16279, 16'd28437};
                15'd5424 : data_rom <= {16'd16282, 16'd28436};
                15'd5425 : data_rom <= {16'd16285, 16'd28434};
                15'd5426 : data_rom <= {16'd16287, 16'd28433};
                15'd5427 : data_rom <= {16'd16290, 16'd28431};
                15'd5428 : data_rom <= {16'd16293, 16'd28430};
                15'd5429 : data_rom <= {16'd16295, 16'd28428};
                15'd5430 : data_rom <= {16'd16298, 16'd28427};
                15'd5431 : data_rom <= {16'd16301, 16'd28425};
                15'd5432 : data_rom <= {16'd16304, 16'd28423};
                15'd5433 : data_rom <= {16'd16306, 16'd28422};
                15'd5434 : data_rom <= {16'd16309, 16'd28420};
                15'd5435 : data_rom <= {16'd16312, 16'd28419};
                15'd5436 : data_rom <= {16'd16315, 16'd28417};
                15'd5437 : data_rom <= {16'd16317, 16'd28416};
                15'd5438 : data_rom <= {16'd16320, 16'd28414};
                15'd5439 : data_rom <= {16'd16323, 16'd28412};
                15'd5440 : data_rom <= {16'd16325, 16'd28411};
                15'd5441 : data_rom <= {16'd16328, 16'd28409};
                15'd5442 : data_rom <= {16'd16331, 16'd28408};
                15'd5443 : data_rom <= {16'd16334, 16'd28406};
                15'd5444 : data_rom <= {16'd16336, 16'd28405};
                15'd5445 : data_rom <= {16'd16339, 16'd28403};
                15'd5446 : data_rom <= {16'd16342, 16'd28401};
                15'd5447 : data_rom <= {16'd16344, 16'd28400};
                15'd5448 : data_rom <= {16'd16347, 16'd28398};
                15'd5449 : data_rom <= {16'd16350, 16'd28397};
                15'd5450 : data_rom <= {16'd16353, 16'd28395};
                15'd5451 : data_rom <= {16'd16355, 16'd28394};
                15'd5452 : data_rom <= {16'd16358, 16'd28392};
                15'd5453 : data_rom <= {16'd16361, 16'd28391};
                15'd5454 : data_rom <= {16'd16364, 16'd28389};
                15'd5455 : data_rom <= {16'd16366, 16'd28387};
                15'd5456 : data_rom <= {16'd16369, 16'd28386};
                15'd5457 : data_rom <= {16'd16372, 16'd28384};
                15'd5458 : data_rom <= {16'd16374, 16'd28383};
                15'd5459 : data_rom <= {16'd16377, 16'd28381};
                15'd5460 : data_rom <= {16'd16380, 16'd28380};
                15'd5461 : data_rom <= {16'd16383, 16'd28378};
                15'd5462 : data_rom <= {16'd16385, 16'd28376};
                15'd5463 : data_rom <= {16'd16388, 16'd28375};
                15'd5464 : data_rom <= {16'd16391, 16'd28373};
                15'd5465 : data_rom <= {16'd16393, 16'd28372};
                15'd5466 : data_rom <= {16'd16396, 16'd28370};
                15'd5467 : data_rom <= {16'd16399, 16'd28369};
                15'd5468 : data_rom <= {16'd16402, 16'd28367};
                15'd5469 : data_rom <= {16'd16404, 16'd28365};
                15'd5470 : data_rom <= {16'd16407, 16'd28364};
                15'd5471 : data_rom <= {16'd16410, 16'd28362};
                15'd5472 : data_rom <= {16'd16412, 16'd28361};
                15'd5473 : data_rom <= {16'd16415, 16'd28359};
                15'd5474 : data_rom <= {16'd16418, 16'd28358};
                15'd5475 : data_rom <= {16'd16421, 16'd28356};
                15'd5476 : data_rom <= {16'd16423, 16'd28354};
                15'd5477 : data_rom <= {16'd16426, 16'd28353};
                15'd5478 : data_rom <= {16'd16429, 16'd28351};
                15'd5479 : data_rom <= {16'd16432, 16'd28350};
                15'd5480 : data_rom <= {16'd16434, 16'd28348};
                15'd5481 : data_rom <= {16'd16437, 16'd28346};
                15'd5482 : data_rom <= {16'd16440, 16'd28345};
                15'd5483 : data_rom <= {16'd16442, 16'd28343};
                15'd5484 : data_rom <= {16'd16445, 16'd28342};
                15'd5485 : data_rom <= {16'd16448, 16'd28340};
                15'd5486 : data_rom <= {16'd16451, 16'd28339};
                15'd5487 : data_rom <= {16'd16453, 16'd28337};
                15'd5488 : data_rom <= {16'd16456, 16'd28335};
                15'd5489 : data_rom <= {16'd16459, 16'd28334};
                15'd5490 : data_rom <= {16'd16461, 16'd28332};
                15'd5491 : data_rom <= {16'd16464, 16'd28331};
                15'd5492 : data_rom <= {16'd16467, 16'd28329};
                15'd5493 : data_rom <= {16'd16470, 16'd28328};
                15'd5494 : data_rom <= {16'd16472, 16'd28326};
                15'd5495 : data_rom <= {16'd16475, 16'd28324};
                15'd5496 : data_rom <= {16'd16478, 16'd28323};
                15'd5497 : data_rom <= {16'd16480, 16'd28321};
                15'd5498 : data_rom <= {16'd16483, 16'd28320};
                15'd5499 : data_rom <= {16'd16486, 16'd28318};
                15'd5500 : data_rom <= {16'd16489, 16'd28316};
                15'd5501 : data_rom <= {16'd16491, 16'd28315};
                15'd5502 : data_rom <= {16'd16494, 16'd28313};
                15'd5503 : data_rom <= {16'd16497, 16'd28312};
                15'd5504 : data_rom <= {16'd16499, 16'd28310};
                15'd5505 : data_rom <= {16'd16502, 16'd28309};
                15'd5506 : data_rom <= {16'd16505, 16'd28307};
                15'd5507 : data_rom <= {16'd16508, 16'd28305};
                15'd5508 : data_rom <= {16'd16510, 16'd28304};
                15'd5509 : data_rom <= {16'd16513, 16'd28302};
                15'd5510 : data_rom <= {16'd16516, 16'd28301};
                15'd5511 : data_rom <= {16'd16518, 16'd28299};
                15'd5512 : data_rom <= {16'd16521, 16'd28298};
                15'd5513 : data_rom <= {16'd16524, 16'd28296};
                15'd5514 : data_rom <= {16'd16527, 16'd28294};
                15'd5515 : data_rom <= {16'd16529, 16'd28293};
                15'd5516 : data_rom <= {16'd16532, 16'd28291};
                15'd5517 : data_rom <= {16'd16535, 16'd28290};
                15'd5518 : data_rom <= {16'd16537, 16'd28288};
                15'd5519 : data_rom <= {16'd16540, 16'd28286};
                15'd5520 : data_rom <= {16'd16543, 16'd28285};
                15'd5521 : data_rom <= {16'd16546, 16'd28283};
                15'd5522 : data_rom <= {16'd16548, 16'd28282};
                15'd5523 : data_rom <= {16'd16551, 16'd28280};
                15'd5524 : data_rom <= {16'd16554, 16'd28278};
                15'd5525 : data_rom <= {16'd16556, 16'd28277};
                15'd5526 : data_rom <= {16'd16559, 16'd28275};
                15'd5527 : data_rom <= {16'd16562, 16'd28274};
                15'd5528 : data_rom <= {16'd16565, 16'd28272};
                15'd5529 : data_rom <= {16'd16567, 16'd28271};
                15'd5530 : data_rom <= {16'd16570, 16'd28269};
                15'd5531 : data_rom <= {16'd16573, 16'd28267};
                15'd5532 : data_rom <= {16'd16575, 16'd28266};
                15'd5533 : data_rom <= {16'd16578, 16'd28264};
                15'd5534 : data_rom <= {16'd16581, 16'd28263};
                15'd5535 : data_rom <= {16'd16584, 16'd28261};
                15'd5536 : data_rom <= {16'd16586, 16'd28259};
                15'd5537 : data_rom <= {16'd16589, 16'd28258};
                15'd5538 : data_rom <= {16'd16592, 16'd28256};
                15'd5539 : data_rom <= {16'd16594, 16'd28255};
                15'd5540 : data_rom <= {16'd16597, 16'd28253};
                15'd5541 : data_rom <= {16'd16600, 16'd28251};
                15'd5542 : data_rom <= {16'd16602, 16'd28250};
                15'd5543 : data_rom <= {16'd16605, 16'd28248};
                15'd5544 : data_rom <= {16'd16608, 16'd28247};
                15'd5545 : data_rom <= {16'd16611, 16'd28245};
                15'd5546 : data_rom <= {16'd16613, 16'd28244};
                15'd5547 : data_rom <= {16'd16616, 16'd28242};
                15'd5548 : data_rom <= {16'd16619, 16'd28240};
                15'd5549 : data_rom <= {16'd16621, 16'd28239};
                15'd5550 : data_rom <= {16'd16624, 16'd28237};
                15'd5551 : data_rom <= {16'd16627, 16'd28236};
                15'd5552 : data_rom <= {16'd16630, 16'd28234};
                15'd5553 : data_rom <= {16'd16632, 16'd28232};
                15'd5554 : data_rom <= {16'd16635, 16'd28231};
                15'd5555 : data_rom <= {16'd16638, 16'd28229};
                15'd5556 : data_rom <= {16'd16640, 16'd28228};
                15'd5557 : data_rom <= {16'd16643, 16'd28226};
                15'd5558 : data_rom <= {16'd16646, 16'd28224};
                15'd5559 : data_rom <= {16'd16648, 16'd28223};
                15'd5560 : data_rom <= {16'd16651, 16'd28221};
                15'd5561 : data_rom <= {16'd16654, 16'd28220};
                15'd5562 : data_rom <= {16'd16657, 16'd28218};
                15'd5563 : data_rom <= {16'd16659, 16'd28216};
                15'd5564 : data_rom <= {16'd16662, 16'd28215};
                15'd5565 : data_rom <= {16'd16665, 16'd28213};
                15'd5566 : data_rom <= {16'd16667, 16'd28212};
                15'd5567 : data_rom <= {16'd16670, 16'd28210};
                15'd5568 : data_rom <= {16'd16673, 16'd28208};
                15'd5569 : data_rom <= {16'd16676, 16'd28207};
                15'd5570 : data_rom <= {16'd16678, 16'd28205};
                15'd5571 : data_rom <= {16'd16681, 16'd28204};
                15'd5572 : data_rom <= {16'd16684, 16'd28202};
                15'd5573 : data_rom <= {16'd16686, 16'd28200};
                15'd5574 : data_rom <= {16'd16689, 16'd28199};
                15'd5575 : data_rom <= {16'd16692, 16'd28197};
                15'd5576 : data_rom <= {16'd16694, 16'd28196};
                15'd5577 : data_rom <= {16'd16697, 16'd28194};
                15'd5578 : data_rom <= {16'd16700, 16'd28192};
                15'd5579 : data_rom <= {16'd16703, 16'd28191};
                15'd5580 : data_rom <= {16'd16705, 16'd28189};
                15'd5581 : data_rom <= {16'd16708, 16'd28188};
                15'd5582 : data_rom <= {16'd16711, 16'd28186};
                15'd5583 : data_rom <= {16'd16713, 16'd28184};
                15'd5584 : data_rom <= {16'd16716, 16'd28183};
                15'd5585 : data_rom <= {16'd16719, 16'd28181};
                15'd5586 : data_rom <= {16'd16721, 16'd28180};
                15'd5587 : data_rom <= {16'd16724, 16'd28178};
                15'd5588 : data_rom <= {16'd16727, 16'd28176};
                15'd5589 : data_rom <= {16'd16730, 16'd28175};
                15'd5590 : data_rom <= {16'd16732, 16'd28173};
                15'd5591 : data_rom <= {16'd16735, 16'd28172};
                15'd5592 : data_rom <= {16'd16738, 16'd28170};
                15'd5593 : data_rom <= {16'd16740, 16'd28168};
                15'd5594 : data_rom <= {16'd16743, 16'd28167};
                15'd5595 : data_rom <= {16'd16746, 16'd28165};
                15'd5596 : data_rom <= {16'd16748, 16'd28164};
                15'd5597 : data_rom <= {16'd16751, 16'd28162};
                15'd5598 : data_rom <= {16'd16754, 16'd28160};
                15'd5599 : data_rom <= {16'd16757, 16'd28159};
                15'd5600 : data_rom <= {16'd16759, 16'd28157};
                15'd5601 : data_rom <= {16'd16762, 16'd28156};
                15'd5602 : data_rom <= {16'd16765, 16'd28154};
                15'd5603 : data_rom <= {16'd16767, 16'd28152};
                15'd5604 : data_rom <= {16'd16770, 16'd28151};
                15'd5605 : data_rom <= {16'd16773, 16'd28149};
                15'd5606 : data_rom <= {16'd16775, 16'd28147};
                15'd5607 : data_rom <= {16'd16778, 16'd28146};
                15'd5608 : data_rom <= {16'd16781, 16'd28144};
                15'd5609 : data_rom <= {16'd16784, 16'd28143};
                15'd5610 : data_rom <= {16'd16786, 16'd28141};
                15'd5611 : data_rom <= {16'd16789, 16'd28139};
                15'd5612 : data_rom <= {16'd16792, 16'd28138};
                15'd5613 : data_rom <= {16'd16794, 16'd28136};
                15'd5614 : data_rom <= {16'd16797, 16'd28135};
                15'd5615 : data_rom <= {16'd16800, 16'd28133};
                15'd5616 : data_rom <= {16'd16802, 16'd28131};
                15'd5617 : data_rom <= {16'd16805, 16'd28130};
                15'd5618 : data_rom <= {16'd16808, 16'd28128};
                15'd5619 : data_rom <= {16'd16811, 16'd28127};
                15'd5620 : data_rom <= {16'd16813, 16'd28125};
                15'd5621 : data_rom <= {16'd16816, 16'd28123};
                15'd5622 : data_rom <= {16'd16819, 16'd28122};
                15'd5623 : data_rom <= {16'd16821, 16'd28120};
                15'd5624 : data_rom <= {16'd16824, 16'd28118};
                15'd5625 : data_rom <= {16'd16827, 16'd28117};
                15'd5626 : data_rom <= {16'd16829, 16'd28115};
                15'd5627 : data_rom <= {16'd16832, 16'd28114};
                15'd5628 : data_rom <= {16'd16835, 16'd28112};
                15'd5629 : data_rom <= {16'd16838, 16'd28110};
                15'd5630 : data_rom <= {16'd16840, 16'd28109};
                15'd5631 : data_rom <= {16'd16843, 16'd28107};
                15'd5632 : data_rom <= {16'd16846, 16'd28106};
                15'd5633 : data_rom <= {16'd16848, 16'd28104};
                15'd5634 : data_rom <= {16'd16851, 16'd28102};
                15'd5635 : data_rom <= {16'd16854, 16'd28101};
                15'd5636 : data_rom <= {16'd16856, 16'd28099};
                15'd5637 : data_rom <= {16'd16859, 16'd28097};
                15'd5638 : data_rom <= {16'd16862, 16'd28096};
                15'd5639 : data_rom <= {16'd16864, 16'd28094};
                15'd5640 : data_rom <= {16'd16867, 16'd28093};
                15'd5641 : data_rom <= {16'd16870, 16'd28091};
                15'd5642 : data_rom <= {16'd16873, 16'd28089};
                15'd5643 : data_rom <= {16'd16875, 16'd28088};
                15'd5644 : data_rom <= {16'd16878, 16'd28086};
                15'd5645 : data_rom <= {16'd16881, 16'd28085};
                15'd5646 : data_rom <= {16'd16883, 16'd28083};
                15'd5647 : data_rom <= {16'd16886, 16'd28081};
                15'd5648 : data_rom <= {16'd16889, 16'd28080};
                15'd5649 : data_rom <= {16'd16891, 16'd28078};
                15'd5650 : data_rom <= {16'd16894, 16'd28076};
                15'd5651 : data_rom <= {16'd16897, 16'd28075};
                15'd5652 : data_rom <= {16'd16899, 16'd28073};
                15'd5653 : data_rom <= {16'd16902, 16'd28072};
                15'd5654 : data_rom <= {16'd16905, 16'd28070};
                15'd5655 : data_rom <= {16'd16908, 16'd28068};
                15'd5656 : data_rom <= {16'd16910, 16'd28067};
                15'd5657 : data_rom <= {16'd16913, 16'd28065};
                15'd5658 : data_rom <= {16'd16916, 16'd28063};
                15'd5659 : data_rom <= {16'd16918, 16'd28062};
                15'd5660 : data_rom <= {16'd16921, 16'd28060};
                15'd5661 : data_rom <= {16'd16924, 16'd28059};
                15'd5662 : data_rom <= {16'd16926, 16'd28057};
                15'd5663 : data_rom <= {16'd16929, 16'd28055};
                15'd5664 : data_rom <= {16'd16932, 16'd28054};
                15'd5665 : data_rom <= {16'd16934, 16'd28052};
                15'd5666 : data_rom <= {16'd16937, 16'd28050};
                15'd5667 : data_rom <= {16'd16940, 16'd28049};
                15'd5668 : data_rom <= {16'd16943, 16'd28047};
                15'd5669 : data_rom <= {16'd16945, 16'd28046};
                15'd5670 : data_rom <= {16'd16948, 16'd28044};
                15'd5671 : data_rom <= {16'd16951, 16'd28042};
                15'd5672 : data_rom <= {16'd16953, 16'd28041};
                15'd5673 : data_rom <= {16'd16956, 16'd28039};
                15'd5674 : data_rom <= {16'd16959, 16'd28037};
                15'd5675 : data_rom <= {16'd16961, 16'd28036};
                15'd5676 : data_rom <= {16'd16964, 16'd28034};
                15'd5677 : data_rom <= {16'd16967, 16'd28033};
                15'd5678 : data_rom <= {16'd16969, 16'd28031};
                15'd5679 : data_rom <= {16'd16972, 16'd28029};
                15'd5680 : data_rom <= {16'd16975, 16'd28028};
                15'd5681 : data_rom <= {16'd16977, 16'd28026};
                15'd5682 : data_rom <= {16'd16980, 16'd28024};
                15'd5683 : data_rom <= {16'd16983, 16'd28023};
                15'd5684 : data_rom <= {16'd16986, 16'd28021};
                15'd5685 : data_rom <= {16'd16988, 16'd28020};
                15'd5686 : data_rom <= {16'd16991, 16'd28018};
                15'd5687 : data_rom <= {16'd16994, 16'd28016};
                15'd5688 : data_rom <= {16'd16996, 16'd28015};
                15'd5689 : data_rom <= {16'd16999, 16'd28013};
                15'd5690 : data_rom <= {16'd17002, 16'd28011};
                15'd5691 : data_rom <= {16'd17004, 16'd28010};
                15'd5692 : data_rom <= {16'd17007, 16'd28008};
                15'd5693 : data_rom <= {16'd17010, 16'd28007};
                15'd5694 : data_rom <= {16'd17012, 16'd28005};
                15'd5695 : data_rom <= {16'd17015, 16'd28003};
                15'd5696 : data_rom <= {16'd17018, 16'd28002};
                15'd5697 : data_rom <= {16'd17020, 16'd28000};
                15'd5698 : data_rom <= {16'd17023, 16'd27998};
                15'd5699 : data_rom <= {16'd17026, 16'd27997};
                15'd5700 : data_rom <= {16'd17028, 16'd27995};
                15'd5701 : data_rom <= {16'd17031, 16'd27994};
                15'd5702 : data_rom <= {16'd17034, 16'd27992};
                15'd5703 : data_rom <= {16'd17037, 16'd27990};
                15'd5704 : data_rom <= {16'd17039, 16'd27989};
                15'd5705 : data_rom <= {16'd17042, 16'd27987};
                15'd5706 : data_rom <= {16'd17045, 16'd27985};
                15'd5707 : data_rom <= {16'd17047, 16'd27984};
                15'd5708 : data_rom <= {16'd17050, 16'd27982};
                15'd5709 : data_rom <= {16'd17053, 16'd27980};
                15'd5710 : data_rom <= {16'd17055, 16'd27979};
                15'd5711 : data_rom <= {16'd17058, 16'd27977};
                15'd5712 : data_rom <= {16'd17061, 16'd27976};
                15'd5713 : data_rom <= {16'd17063, 16'd27974};
                15'd5714 : data_rom <= {16'd17066, 16'd27972};
                15'd5715 : data_rom <= {16'd17069, 16'd27971};
                15'd5716 : data_rom <= {16'd17071, 16'd27969};
                15'd5717 : data_rom <= {16'd17074, 16'd27967};
                15'd5718 : data_rom <= {16'd17077, 16'd27966};
                15'd5719 : data_rom <= {16'd17079, 16'd27964};
                15'd5720 : data_rom <= {16'd17082, 16'd27962};
                15'd5721 : data_rom <= {16'd17085, 16'd27961};
                15'd5722 : data_rom <= {16'd17087, 16'd27959};
                15'd5723 : data_rom <= {16'd17090, 16'd27958};
                15'd5724 : data_rom <= {16'd17093, 16'd27956};
                15'd5725 : data_rom <= {16'd17096, 16'd27954};
                15'd5726 : data_rom <= {16'd17098, 16'd27953};
                15'd5727 : data_rom <= {16'd17101, 16'd27951};
                15'd5728 : data_rom <= {16'd17104, 16'd27949};
                15'd5729 : data_rom <= {16'd17106, 16'd27948};
                15'd5730 : data_rom <= {16'd17109, 16'd27946};
                15'd5731 : data_rom <= {16'd17112, 16'd27944};
                15'd5732 : data_rom <= {16'd17114, 16'd27943};
                15'd5733 : data_rom <= {16'd17117, 16'd27941};
                15'd5734 : data_rom <= {16'd17120, 16'd27939};
                15'd5735 : data_rom <= {16'd17122, 16'd27938};
                15'd5736 : data_rom <= {16'd17125, 16'd27936};
                15'd5737 : data_rom <= {16'd17128, 16'd27935};
                15'd5738 : data_rom <= {16'd17130, 16'd27933};
                15'd5739 : data_rom <= {16'd17133, 16'd27931};
                15'd5740 : data_rom <= {16'd17136, 16'd27930};
                15'd5741 : data_rom <= {16'd17138, 16'd27928};
                15'd5742 : data_rom <= {16'd17141, 16'd27926};
                15'd5743 : data_rom <= {16'd17144, 16'd27925};
                15'd5744 : data_rom <= {16'd17146, 16'd27923};
                15'd5745 : data_rom <= {16'd17149, 16'd27921};
                15'd5746 : data_rom <= {16'd17152, 16'd27920};
                15'd5747 : data_rom <= {16'd17154, 16'd27918};
                15'd5748 : data_rom <= {16'd17157, 16'd27916};
                15'd5749 : data_rom <= {16'd17160, 16'd27915};
                15'd5750 : data_rom <= {16'd17162, 16'd27913};
                15'd5751 : data_rom <= {16'd17165, 16'd27912};
                15'd5752 : data_rom <= {16'd17168, 16'd27910};
                15'd5753 : data_rom <= {16'd17171, 16'd27908};
                15'd5754 : data_rom <= {16'd17173, 16'd27907};
                15'd5755 : data_rom <= {16'd17176, 16'd27905};
                15'd5756 : data_rom <= {16'd17179, 16'd27903};
                15'd5757 : data_rom <= {16'd17181, 16'd27902};
                15'd5758 : data_rom <= {16'd17184, 16'd27900};
                15'd5759 : data_rom <= {16'd17187, 16'd27898};
                15'd5760 : data_rom <= {16'd17189, 16'd27897};
                15'd5761 : data_rom <= {16'd17192, 16'd27895};
                15'd5762 : data_rom <= {16'd17195, 16'd27893};
                15'd5763 : data_rom <= {16'd17197, 16'd27892};
                15'd5764 : data_rom <= {16'd17200, 16'd27890};
                15'd5765 : data_rom <= {16'd17203, 16'd27888};
                15'd5766 : data_rom <= {16'd17205, 16'd27887};
                15'd5767 : data_rom <= {16'd17208, 16'd27885};
                15'd5768 : data_rom <= {16'd17211, 16'd27884};
                15'd5769 : data_rom <= {16'd17213, 16'd27882};
                15'd5770 : data_rom <= {16'd17216, 16'd27880};
                15'd5771 : data_rom <= {16'd17219, 16'd27879};
                15'd5772 : data_rom <= {16'd17221, 16'd27877};
                15'd5773 : data_rom <= {16'd17224, 16'd27875};
                15'd5774 : data_rom <= {16'd17227, 16'd27874};
                15'd5775 : data_rom <= {16'd17229, 16'd27872};
                15'd5776 : data_rom <= {16'd17232, 16'd27870};
                15'd5777 : data_rom <= {16'd17235, 16'd27869};
                15'd5778 : data_rom <= {16'd17237, 16'd27867};
                15'd5779 : data_rom <= {16'd17240, 16'd27865};
                15'd5780 : data_rom <= {16'd17243, 16'd27864};
                15'd5781 : data_rom <= {16'd17245, 16'd27862};
                15'd5782 : data_rom <= {16'd17248, 16'd27860};
                15'd5783 : data_rom <= {16'd17251, 16'd27859};
                15'd5784 : data_rom <= {16'd17253, 16'd27857};
                15'd5785 : data_rom <= {16'd17256, 16'd27855};
                15'd5786 : data_rom <= {16'd17259, 16'd27854};
                15'd5787 : data_rom <= {16'd17261, 16'd27852};
                15'd5788 : data_rom <= {16'd17264, 16'd27850};
                15'd5789 : data_rom <= {16'd17267, 16'd27849};
                15'd5790 : data_rom <= {16'd17269, 16'd27847};
                15'd5791 : data_rom <= {16'd17272, 16'd27846};
                15'd5792 : data_rom <= {16'd17275, 16'd27844};
                15'd5793 : data_rom <= {16'd17277, 16'd27842};
                15'd5794 : data_rom <= {16'd17280, 16'd27841};
                15'd5795 : data_rom <= {16'd17283, 16'd27839};
                15'd5796 : data_rom <= {16'd17285, 16'd27837};
                15'd5797 : data_rom <= {16'd17288, 16'd27836};
                15'd5798 : data_rom <= {16'd17291, 16'd27834};
                15'd5799 : data_rom <= {16'd17293, 16'd27832};
                15'd5800 : data_rom <= {16'd17296, 16'd27831};
                15'd5801 : data_rom <= {16'd17299, 16'd27829};
                15'd5802 : data_rom <= {16'd17301, 16'd27827};
                15'd5803 : data_rom <= {16'd17304, 16'd27826};
                15'd5804 : data_rom <= {16'd17307, 16'd27824};
                15'd5805 : data_rom <= {16'd17309, 16'd27822};
                15'd5806 : data_rom <= {16'd17312, 16'd27821};
                15'd5807 : data_rom <= {16'd17315, 16'd27819};
                15'd5808 : data_rom <= {16'd17317, 16'd27817};
                15'd5809 : data_rom <= {16'd17320, 16'd27816};
                15'd5810 : data_rom <= {16'd17323, 16'd27814};
                15'd5811 : data_rom <= {16'd17325, 16'd27812};
                15'd5812 : data_rom <= {16'd17328, 16'd27811};
                15'd5813 : data_rom <= {16'd17331, 16'd27809};
                15'd5814 : data_rom <= {16'd17333, 16'd27807};
                15'd5815 : data_rom <= {16'd17336, 16'd27806};
                15'd5816 : data_rom <= {16'd17339, 16'd27804};
                15'd5817 : data_rom <= {16'd17341, 16'd27802};
                15'd5818 : data_rom <= {16'd17344, 16'd27801};
                15'd5819 : data_rom <= {16'd17347, 16'd27799};
                15'd5820 : data_rom <= {16'd17349, 16'd27797};
                15'd5821 : data_rom <= {16'd17352, 16'd27796};
                15'd5822 : data_rom <= {16'd17355, 16'd27794};
                15'd5823 : data_rom <= {16'd17357, 16'd27792};
                15'd5824 : data_rom <= {16'd17360, 16'd27791};
                15'd5825 : data_rom <= {16'd17363, 16'd27789};
                15'd5826 : data_rom <= {16'd17365, 16'd27787};
                15'd5827 : data_rom <= {16'd17368, 16'd27786};
                15'd5828 : data_rom <= {16'd17371, 16'd27784};
                15'd5829 : data_rom <= {16'd17373, 16'd27782};
                15'd5830 : data_rom <= {16'd17376, 16'd27781};
                15'd5831 : data_rom <= {16'd17379, 16'd27779};
                15'd5832 : data_rom <= {16'd17381, 16'd27777};
                15'd5833 : data_rom <= {16'd17384, 16'd27776};
                15'd5834 : data_rom <= {16'd17387, 16'd27774};
                15'd5835 : data_rom <= {16'd17389, 16'd27772};
                15'd5836 : data_rom <= {16'd17392, 16'd27771};
                15'd5837 : data_rom <= {16'd17395, 16'd27769};
                15'd5838 : data_rom <= {16'd17397, 16'd27767};
                15'd5839 : data_rom <= {16'd17400, 16'd27766};
                15'd5840 : data_rom <= {16'd17403, 16'd27764};
                15'd5841 : data_rom <= {16'd17405, 16'd27762};
                15'd5842 : data_rom <= {16'd17408, 16'd27761};
                15'd5843 : data_rom <= {16'd17411, 16'd27759};
                15'd5844 : data_rom <= {16'd17413, 16'd27757};
                15'd5845 : data_rom <= {16'd17416, 16'd27756};
                15'd5846 : data_rom <= {16'd17419, 16'd27754};
                15'd5847 : data_rom <= {16'd17421, 16'd27752};
                15'd5848 : data_rom <= {16'd17424, 16'd27751};
                15'd5849 : data_rom <= {16'd17427, 16'd27749};
                15'd5850 : data_rom <= {16'd17429, 16'd27747};
                15'd5851 : data_rom <= {16'd17432, 16'd27746};
                15'd5852 : data_rom <= {16'd17435, 16'd27744};
                15'd5853 : data_rom <= {16'd17437, 16'd27742};
                15'd5854 : data_rom <= {16'd17440, 16'd27741};
                15'd5855 : data_rom <= {16'd17443, 16'd27739};
                15'd5856 : data_rom <= {16'd17445, 16'd27737};
                15'd5857 : data_rom <= {16'd17448, 16'd27736};
                15'd5858 : data_rom <= {16'd17451, 16'd27734};
                15'd5859 : data_rom <= {16'd17453, 16'd27732};
                15'd5860 : data_rom <= {16'd17456, 16'd27731};
                15'd5861 : data_rom <= {16'd17459, 16'd27729};
                15'd5862 : data_rom <= {16'd17461, 16'd27727};
                15'd5863 : data_rom <= {16'd17464, 16'd27726};
                15'd5864 : data_rom <= {16'd17467, 16'd27724};
                15'd5865 : data_rom <= {16'd17469, 16'd27722};
                15'd5866 : data_rom <= {16'd17472, 16'd27721};
                15'd5867 : data_rom <= {16'd17475, 16'd27719};
                15'd5868 : data_rom <= {16'd17477, 16'd27717};
                15'd5869 : data_rom <= {16'd17480, 16'd27716};
                15'd5870 : data_rom <= {16'd17482, 16'd27714};
                15'd5871 : data_rom <= {16'd17485, 16'd27712};
                15'd5872 : data_rom <= {16'd17488, 16'd27711};
                15'd5873 : data_rom <= {16'd17490, 16'd27709};
                15'd5874 : data_rom <= {16'd17493, 16'd27707};
                15'd5875 : data_rom <= {16'd17496, 16'd27705};
                15'd5876 : data_rom <= {16'd17498, 16'd27704};
                15'd5877 : data_rom <= {16'd17501, 16'd27702};
                15'd5878 : data_rom <= {16'd17504, 16'd27700};
                15'd5879 : data_rom <= {16'd17506, 16'd27699};
                15'd5880 : data_rom <= {16'd17509, 16'd27697};
                15'd5881 : data_rom <= {16'd17512, 16'd27695};
                15'd5882 : data_rom <= {16'd17514, 16'd27694};
                15'd5883 : data_rom <= {16'd17517, 16'd27692};
                15'd5884 : data_rom <= {16'd17520, 16'd27690};
                15'd5885 : data_rom <= {16'd17522, 16'd27689};
                15'd5886 : data_rom <= {16'd17525, 16'd27687};
                15'd5887 : data_rom <= {16'd17528, 16'd27685};
                15'd5888 : data_rom <= {16'd17530, 16'd27684};
                15'd5889 : data_rom <= {16'd17533, 16'd27682};
                15'd5890 : data_rom <= {16'd17536, 16'd27680};
                15'd5891 : data_rom <= {16'd17538, 16'd27679};
                15'd5892 : data_rom <= {16'd17541, 16'd27677};
                15'd5893 : data_rom <= {16'd17544, 16'd27675};
                15'd5894 : data_rom <= {16'd17546, 16'd27674};
                15'd5895 : data_rom <= {16'd17549, 16'd27672};
                15'd5896 : data_rom <= {16'd17552, 16'd27670};
                15'd5897 : data_rom <= {16'd17554, 16'd27669};
                15'd5898 : data_rom <= {16'd17557, 16'd27667};
                15'd5899 : data_rom <= {16'd17559, 16'd27665};
                15'd5900 : data_rom <= {16'd17562, 16'd27663};
                15'd5901 : data_rom <= {16'd17565, 16'd27662};
                15'd5902 : data_rom <= {16'd17567, 16'd27660};
                15'd5903 : data_rom <= {16'd17570, 16'd27658};
                15'd5904 : data_rom <= {16'd17573, 16'd27657};
                15'd5905 : data_rom <= {16'd17575, 16'd27655};
                15'd5906 : data_rom <= {16'd17578, 16'd27653};
                15'd5907 : data_rom <= {16'd17581, 16'd27652};
                15'd5908 : data_rom <= {16'd17583, 16'd27650};
                15'd5909 : data_rom <= {16'd17586, 16'd27648};
                15'd5910 : data_rom <= {16'd17589, 16'd27647};
                15'd5911 : data_rom <= {16'd17591, 16'd27645};
                15'd5912 : data_rom <= {16'd17594, 16'd27643};
                15'd5913 : data_rom <= {16'd17597, 16'd27642};
                15'd5914 : data_rom <= {16'd17599, 16'd27640};
                15'd5915 : data_rom <= {16'd17602, 16'd27638};
                15'd5916 : data_rom <= {16'd17605, 16'd27637};
                15'd5917 : data_rom <= {16'd17607, 16'd27635};
                15'd5918 : data_rom <= {16'd17610, 16'd27633};
                15'd5919 : data_rom <= {16'd17612, 16'd27631};
                15'd5920 : data_rom <= {16'd17615, 16'd27630};
                15'd5921 : data_rom <= {16'd17618, 16'd27628};
                15'd5922 : data_rom <= {16'd17620, 16'd27626};
                15'd5923 : data_rom <= {16'd17623, 16'd27625};
                15'd5924 : data_rom <= {16'd17626, 16'd27623};
                15'd5925 : data_rom <= {16'd17628, 16'd27621};
                15'd5926 : data_rom <= {16'd17631, 16'd27620};
                15'd5927 : data_rom <= {16'd17634, 16'd27618};
                15'd5928 : data_rom <= {16'd17636, 16'd27616};
                15'd5929 : data_rom <= {16'd17639, 16'd27615};
                15'd5930 : data_rom <= {16'd17642, 16'd27613};
                15'd5931 : data_rom <= {16'd17644, 16'd27611};
                15'd5932 : data_rom <= {16'd17647, 16'd27609};
                15'd5933 : data_rom <= {16'd17650, 16'd27608};
                15'd5934 : data_rom <= {16'd17652, 16'd27606};
                15'd5935 : data_rom <= {16'd17655, 16'd27604};
                15'd5936 : data_rom <= {16'd17658, 16'd27603};
                15'd5937 : data_rom <= {16'd17660, 16'd27601};
                15'd5938 : data_rom <= {16'd17663, 16'd27599};
                15'd5939 : data_rom <= {16'd17665, 16'd27598};
                15'd5940 : data_rom <= {16'd17668, 16'd27596};
                15'd5941 : data_rom <= {16'd17671, 16'd27594};
                15'd5942 : data_rom <= {16'd17673, 16'd27593};
                15'd5943 : data_rom <= {16'd17676, 16'd27591};
                15'd5944 : data_rom <= {16'd17679, 16'd27589};
                15'd5945 : data_rom <= {16'd17681, 16'd27587};
                15'd5946 : data_rom <= {16'd17684, 16'd27586};
                15'd5947 : data_rom <= {16'd17687, 16'd27584};
                15'd5948 : data_rom <= {16'd17689, 16'd27582};
                15'd5949 : data_rom <= {16'd17692, 16'd27581};
                15'd5950 : data_rom <= {16'd17695, 16'd27579};
                15'd5951 : data_rom <= {16'd17697, 16'd27577};
                15'd5952 : data_rom <= {16'd17700, 16'd27576};
                15'd5953 : data_rom <= {16'd17702, 16'd27574};
                15'd5954 : data_rom <= {16'd17705, 16'd27572};
                15'd5955 : data_rom <= {16'd17708, 16'd27570};
                15'd5956 : data_rom <= {16'd17710, 16'd27569};
                15'd5957 : data_rom <= {16'd17713, 16'd27567};
                15'd5958 : data_rom <= {16'd17716, 16'd27565};
                15'd5959 : data_rom <= {16'd17718, 16'd27564};
                15'd5960 : data_rom <= {16'd17721, 16'd27562};
                15'd5961 : data_rom <= {16'd17724, 16'd27560};
                15'd5962 : data_rom <= {16'd17726, 16'd27559};
                15'd5963 : data_rom <= {16'd17729, 16'd27557};
                15'd5964 : data_rom <= {16'd17732, 16'd27555};
                15'd5965 : data_rom <= {16'd17734, 16'd27554};
                15'd5966 : data_rom <= {16'd17737, 16'd27552};
                15'd5967 : data_rom <= {16'd17739, 16'd27550};
                15'd5968 : data_rom <= {16'd17742, 16'd27548};
                15'd5969 : data_rom <= {16'd17745, 16'd27547};
                15'd5970 : data_rom <= {16'd17747, 16'd27545};
                15'd5971 : data_rom <= {16'd17750, 16'd27543};
                15'd5972 : data_rom <= {16'd17753, 16'd27542};
                15'd5973 : data_rom <= {16'd17755, 16'd27540};
                15'd5974 : data_rom <= {16'd17758, 16'd27538};
                15'd5975 : data_rom <= {16'd17761, 16'd27536};
                15'd5976 : data_rom <= {16'd17763, 16'd27535};
                15'd5977 : data_rom <= {16'd17766, 16'd27533};
                15'd5978 : data_rom <= {16'd17769, 16'd27531};
                15'd5979 : data_rom <= {16'd17771, 16'd27530};
                15'd5980 : data_rom <= {16'd17774, 16'd27528};
                15'd5981 : data_rom <= {16'd17776, 16'd27526};
                15'd5982 : data_rom <= {16'd17779, 16'd27525};
                15'd5983 : data_rom <= {16'd17782, 16'd27523};
                15'd5984 : data_rom <= {16'd17784, 16'd27521};
                15'd5985 : data_rom <= {16'd17787, 16'd27519};
                15'd5986 : data_rom <= {16'd17790, 16'd27518};
                15'd5987 : data_rom <= {16'd17792, 16'd27516};
                15'd5988 : data_rom <= {16'd17795, 16'd27514};
                15'd5989 : data_rom <= {16'd17798, 16'd27513};
                15'd5990 : data_rom <= {16'd17800, 16'd27511};
                15'd5991 : data_rom <= {16'd17803, 16'd27509};
                15'd5992 : data_rom <= {16'd17805, 16'd27508};
                15'd5993 : data_rom <= {16'd17808, 16'd27506};
                15'd5994 : data_rom <= {16'd17811, 16'd27504};
                15'd5995 : data_rom <= {16'd17813, 16'd27502};
                15'd5996 : data_rom <= {16'd17816, 16'd27501};
                15'd5997 : data_rom <= {16'd17819, 16'd27499};
                15'd5998 : data_rom <= {16'd17821, 16'd27497};
                15'd5999 : data_rom <= {16'd17824, 16'd27496};
                15'd6000 : data_rom <= {16'd17827, 16'd27494};
                15'd6001 : data_rom <= {16'd17829, 16'd27492};
                15'd6002 : data_rom <= {16'd17832, 16'd27490};
                15'd6003 : data_rom <= {16'd17834, 16'd27489};
                15'd6004 : data_rom <= {16'd17837, 16'd27487};
                15'd6005 : data_rom <= {16'd17840, 16'd27485};
                15'd6006 : data_rom <= {16'd17842, 16'd27484};
                15'd6007 : data_rom <= {16'd17845, 16'd27482};
                15'd6008 : data_rom <= {16'd17848, 16'd27480};
                15'd6009 : data_rom <= {16'd17850, 16'd27478};
                15'd6010 : data_rom <= {16'd17853, 16'd27477};
                15'd6011 : data_rom <= {16'd17856, 16'd27475};
                15'd6012 : data_rom <= {16'd17858, 16'd27473};
                15'd6013 : data_rom <= {16'd17861, 16'd27472};
                15'd6014 : data_rom <= {16'd17863, 16'd27470};
                15'd6015 : data_rom <= {16'd17866, 16'd27468};
                15'd6016 : data_rom <= {16'd17869, 16'd27466};
                15'd6017 : data_rom <= {16'd17871, 16'd27465};
                15'd6018 : data_rom <= {16'd17874, 16'd27463};
                15'd6019 : data_rom <= {16'd17877, 16'd27461};
                15'd6020 : data_rom <= {16'd17879, 16'd27460};
                15'd6021 : data_rom <= {16'd17882, 16'd27458};
                15'd6022 : data_rom <= {16'd17884, 16'd27456};
                15'd6023 : data_rom <= {16'd17887, 16'd27454};
                15'd6024 : data_rom <= {16'd17890, 16'd27453};
                15'd6025 : data_rom <= {16'd17892, 16'd27451};
                15'd6026 : data_rom <= {16'd17895, 16'd27449};
                15'd6027 : data_rom <= {16'd17898, 16'd27448};
                15'd6028 : data_rom <= {16'd17900, 16'd27446};
                15'd6029 : data_rom <= {16'd17903, 16'd27444};
                15'd6030 : data_rom <= {16'd17906, 16'd27442};
                15'd6031 : data_rom <= {16'd17908, 16'd27441};
                15'd6032 : data_rom <= {16'd17911, 16'd27439};
                15'd6033 : data_rom <= {16'd17913, 16'd27437};
                15'd6034 : data_rom <= {16'd17916, 16'd27436};
                15'd6035 : data_rom <= {16'd17919, 16'd27434};
                15'd6036 : data_rom <= {16'd17921, 16'd27432};
                15'd6037 : data_rom <= {16'd17924, 16'd27430};
                15'd6038 : data_rom <= {16'd17927, 16'd27429};
                15'd6039 : data_rom <= {16'd17929, 16'd27427};
                15'd6040 : data_rom <= {16'd17932, 16'd27425};
                15'd6041 : data_rom <= {16'd17934, 16'd27424};
                15'd6042 : data_rom <= {16'd17937, 16'd27422};
                15'd6043 : data_rom <= {16'd17940, 16'd27420};
                15'd6044 : data_rom <= {16'd17942, 16'd27418};
                15'd6045 : data_rom <= {16'd17945, 16'd27417};
                15'd6046 : data_rom <= {16'd17948, 16'd27415};
                15'd6047 : data_rom <= {16'd17950, 16'd27413};
                15'd6048 : data_rom <= {16'd17953, 16'd27412};
                15'd6049 : data_rom <= {16'd17956, 16'd27410};
                15'd6050 : data_rom <= {16'd17958, 16'd27408};
                15'd6051 : data_rom <= {16'd17961, 16'd27406};
                15'd6052 : data_rom <= {16'd17963, 16'd27405};
                15'd6053 : data_rom <= {16'd17966, 16'd27403};
                15'd6054 : data_rom <= {16'd17969, 16'd27401};
                15'd6055 : data_rom <= {16'd17971, 16'd27399};
                15'd6056 : data_rom <= {16'd17974, 16'd27398};
                15'd6057 : data_rom <= {16'd17977, 16'd27396};
                15'd6058 : data_rom <= {16'd17979, 16'd27394};
                15'd6059 : data_rom <= {16'd17982, 16'd27393};
                15'd6060 : data_rom <= {16'd17984, 16'd27391};
                15'd6061 : data_rom <= {16'd17987, 16'd27389};
                15'd6062 : data_rom <= {16'd17990, 16'd27387};
                15'd6063 : data_rom <= {16'd17992, 16'd27386};
                15'd6064 : data_rom <= {16'd17995, 16'd27384};
                15'd6065 : data_rom <= {16'd17998, 16'd27382};
                15'd6066 : data_rom <= {16'd18000, 16'd27380};
                15'd6067 : data_rom <= {16'd18003, 16'd27379};
                15'd6068 : data_rom <= {16'd18005, 16'd27377};
                15'd6069 : data_rom <= {16'd18008, 16'd27375};
                15'd6070 : data_rom <= {16'd18011, 16'd27374};
                15'd6071 : data_rom <= {16'd18013, 16'd27372};
                15'd6072 : data_rom <= {16'd18016, 16'd27370};
                15'd6073 : data_rom <= {16'd18019, 16'd27368};
                15'd6074 : data_rom <= {16'd18021, 16'd27367};
                15'd6075 : data_rom <= {16'd18024, 16'd27365};
                15'd6076 : data_rom <= {16'd18026, 16'd27363};
                15'd6077 : data_rom <= {16'd18029, 16'd27361};
                15'd6078 : data_rom <= {16'd18032, 16'd27360};
                15'd6079 : data_rom <= {16'd18034, 16'd27358};
                15'd6080 : data_rom <= {16'd18037, 16'd27356};
                15'd6081 : data_rom <= {16'd18040, 16'd27355};
                15'd6082 : data_rom <= {16'd18042, 16'd27353};
                15'd6083 : data_rom <= {16'd18045, 16'd27351};
                15'd6084 : data_rom <= {16'd18047, 16'd27349};
                15'd6085 : data_rom <= {16'd18050, 16'd27348};
                15'd6086 : data_rom <= {16'd18053, 16'd27346};
                15'd6087 : data_rom <= {16'd18055, 16'd27344};
                15'd6088 : data_rom <= {16'd18058, 16'd27342};
                15'd6089 : data_rom <= {16'd18060, 16'd27341};
                15'd6090 : data_rom <= {16'd18063, 16'd27339};
                15'd6091 : data_rom <= {16'd18066, 16'd27337};
                15'd6092 : data_rom <= {16'd18068, 16'd27336};
                15'd6093 : data_rom <= {16'd18071, 16'd27334};
                15'd6094 : data_rom <= {16'd18074, 16'd27332};
                15'd6095 : data_rom <= {16'd18076, 16'd27330};
                15'd6096 : data_rom <= {16'd18079, 16'd27329};
                15'd6097 : data_rom <= {16'd18081, 16'd27327};
                15'd6098 : data_rom <= {16'd18084, 16'd27325};
                15'd6099 : data_rom <= {16'd18087, 16'd27323};
                15'd6100 : data_rom <= {16'd18089, 16'd27322};
                15'd6101 : data_rom <= {16'd18092, 16'd27320};
                15'd6102 : data_rom <= {16'd18095, 16'd27318};
                15'd6103 : data_rom <= {16'd18097, 16'd27316};
                15'd6104 : data_rom <= {16'd18100, 16'd27315};
                15'd6105 : data_rom <= {16'd18102, 16'd27313};
                15'd6106 : data_rom <= {16'd18105, 16'd27311};
                15'd6107 : data_rom <= {16'd18108, 16'd27310};
                15'd6108 : data_rom <= {16'd18110, 16'd27308};
                15'd6109 : data_rom <= {16'd18113, 16'd27306};
                15'd6110 : data_rom <= {16'd18116, 16'd27304};
                15'd6111 : data_rom <= {16'd18118, 16'd27303};
                15'd6112 : data_rom <= {16'd18121, 16'd27301};
                15'd6113 : data_rom <= {16'd18123, 16'd27299};
                15'd6114 : data_rom <= {16'd18126, 16'd27297};
                15'd6115 : data_rom <= {16'd18129, 16'd27296};
                15'd6116 : data_rom <= {16'd18131, 16'd27294};
                15'd6117 : data_rom <= {16'd18134, 16'd27292};
                15'd6118 : data_rom <= {16'd18136, 16'd27290};
                15'd6119 : data_rom <= {16'd18139, 16'd27289};
                15'd6120 : data_rom <= {16'd18142, 16'd27287};
                15'd6121 : data_rom <= {16'd18144, 16'd27285};
                15'd6122 : data_rom <= {16'd18147, 16'd27283};
                15'd6123 : data_rom <= {16'd18150, 16'd27282};
                15'd6124 : data_rom <= {16'd18152, 16'd27280};
                15'd6125 : data_rom <= {16'd18155, 16'd27278};
                15'd6126 : data_rom <= {16'd18157, 16'd27276};
                15'd6127 : data_rom <= {16'd18160, 16'd27275};
                15'd6128 : data_rom <= {16'd18163, 16'd27273};
                15'd6129 : data_rom <= {16'd18165, 16'd27271};
                15'd6130 : data_rom <= {16'd18168, 16'd27270};
                15'd6131 : data_rom <= {16'd18170, 16'd27268};
                15'd6132 : data_rom <= {16'd18173, 16'd27266};
                15'd6133 : data_rom <= {16'd18176, 16'd27264};
                15'd6134 : data_rom <= {16'd18178, 16'd27263};
                15'd6135 : data_rom <= {16'd18181, 16'd27261};
                15'd6136 : data_rom <= {16'd18184, 16'd27259};
                15'd6137 : data_rom <= {16'd18186, 16'd27257};
                15'd6138 : data_rom <= {16'd18189, 16'd27256};
                15'd6139 : data_rom <= {16'd18191, 16'd27254};
                15'd6140 : data_rom <= {16'd18194, 16'd27252};
                15'd6141 : data_rom <= {16'd18197, 16'd27250};
                15'd6142 : data_rom <= {16'd18199, 16'd27249};
                15'd6143 : data_rom <= {16'd18202, 16'd27247};
                15'd6144 : data_rom <= {16'd18204, 16'd27245};
                15'd6145 : data_rom <= {16'd18207, 16'd27243};
                15'd6146 : data_rom <= {16'd18210, 16'd27242};
                15'd6147 : data_rom <= {16'd18212, 16'd27240};
                15'd6148 : data_rom <= {16'd18215, 16'd27238};
                15'd6149 : data_rom <= {16'd18217, 16'd27236};
                15'd6150 : data_rom <= {16'd18220, 16'd27235};
                15'd6151 : data_rom <= {16'd18223, 16'd27233};
                15'd6152 : data_rom <= {16'd18225, 16'd27231};
                15'd6153 : data_rom <= {16'd18228, 16'd27229};
                15'd6154 : data_rom <= {16'd18231, 16'd27228};
                15'd6155 : data_rom <= {16'd18233, 16'd27226};
                15'd6156 : data_rom <= {16'd18236, 16'd27224};
                15'd6157 : data_rom <= {16'd18238, 16'd27222};
                15'd6158 : data_rom <= {16'd18241, 16'd27221};
                15'd6159 : data_rom <= {16'd18244, 16'd27219};
                15'd6160 : data_rom <= {16'd18246, 16'd27217};
                15'd6161 : data_rom <= {16'd18249, 16'd27215};
                15'd6162 : data_rom <= {16'd18251, 16'd27214};
                15'd6163 : data_rom <= {16'd18254, 16'd27212};
                15'd6164 : data_rom <= {16'd18257, 16'd27210};
                15'd6165 : data_rom <= {16'd18259, 16'd27208};
                15'd6166 : data_rom <= {16'd18262, 16'd27207};
                15'd6167 : data_rom <= {16'd18264, 16'd27205};
                15'd6168 : data_rom <= {16'd18267, 16'd27203};
                15'd6169 : data_rom <= {16'd18270, 16'd27201};
                15'd6170 : data_rom <= {16'd18272, 16'd27200};
                15'd6171 : data_rom <= {16'd18275, 16'd27198};
                15'd6172 : data_rom <= {16'd18277, 16'd27196};
                15'd6173 : data_rom <= {16'd18280, 16'd27194};
                15'd6174 : data_rom <= {16'd18283, 16'd27193};
                15'd6175 : data_rom <= {16'd18285, 16'd27191};
                15'd6176 : data_rom <= {16'd18288, 16'd27189};
                15'd6177 : data_rom <= {16'd18291, 16'd27187};
                15'd6178 : data_rom <= {16'd18293, 16'd27186};
                15'd6179 : data_rom <= {16'd18296, 16'd27184};
                15'd6180 : data_rom <= {16'd18298, 16'd27182};
                15'd6181 : data_rom <= {16'd18301, 16'd27180};
                15'd6182 : data_rom <= {16'd18304, 16'd27179};
                15'd6183 : data_rom <= {16'd18306, 16'd27177};
                15'd6184 : data_rom <= {16'd18309, 16'd27175};
                15'd6185 : data_rom <= {16'd18311, 16'd27173};
                15'd6186 : data_rom <= {16'd18314, 16'd27172};
                15'd6187 : data_rom <= {16'd18317, 16'd27170};
                15'd6188 : data_rom <= {16'd18319, 16'd27168};
                15'd6189 : data_rom <= {16'd18322, 16'd27166};
                15'd6190 : data_rom <= {16'd18324, 16'd27165};
                15'd6191 : data_rom <= {16'd18327, 16'd27163};
                15'd6192 : data_rom <= {16'd18330, 16'd27161};
                15'd6193 : data_rom <= {16'd18332, 16'd27159};
                15'd6194 : data_rom <= {16'd18335, 16'd27158};
                15'd6195 : data_rom <= {16'd18337, 16'd27156};
                15'd6196 : data_rom <= {16'd18340, 16'd27154};
                15'd6197 : data_rom <= {16'd18343, 16'd27152};
                15'd6198 : data_rom <= {16'd18345, 16'd27150};
                15'd6199 : data_rom <= {16'd18348, 16'd27149};
                15'd6200 : data_rom <= {16'd18350, 16'd27147};
                15'd6201 : data_rom <= {16'd18353, 16'd27145};
                15'd6202 : data_rom <= {16'd18356, 16'd27143};
                15'd6203 : data_rom <= {16'd18358, 16'd27142};
                15'd6204 : data_rom <= {16'd18361, 16'd27140};
                15'd6205 : data_rom <= {16'd18363, 16'd27138};
                15'd6206 : data_rom <= {16'd18366, 16'd27136};
                15'd6207 : data_rom <= {16'd18369, 16'd27135};
                15'd6208 : data_rom <= {16'd18371, 16'd27133};
                15'd6209 : data_rom <= {16'd18374, 16'd27131};
                15'd6210 : data_rom <= {16'd18376, 16'd27129};
                15'd6211 : data_rom <= {16'd18379, 16'd27128};
                15'd6212 : data_rom <= {16'd18382, 16'd27126};
                15'd6213 : data_rom <= {16'd18384, 16'd27124};
                15'd6214 : data_rom <= {16'd18387, 16'd27122};
                15'd6215 : data_rom <= {16'd18389, 16'd27121};
                15'd6216 : data_rom <= {16'd18392, 16'd27119};
                15'd6217 : data_rom <= {16'd18395, 16'd27117};
                15'd6218 : data_rom <= {16'd18397, 16'd27115};
                15'd6219 : data_rom <= {16'd18400, 16'd27114};
                15'd6220 : data_rom <= {16'd18402, 16'd27112};
                15'd6221 : data_rom <= {16'd18405, 16'd27110};
                15'd6222 : data_rom <= {16'd18408, 16'd27108};
                15'd6223 : data_rom <= {16'd18410, 16'd27106};
                15'd6224 : data_rom <= {16'd18413, 16'd27105};
                15'd6225 : data_rom <= {16'd18415, 16'd27103};
                15'd6226 : data_rom <= {16'd18418, 16'd27101};
                15'd6227 : data_rom <= {16'd18421, 16'd27099};
                15'd6228 : data_rom <= {16'd18423, 16'd27098};
                15'd6229 : data_rom <= {16'd18426, 16'd27096};
                15'd6230 : data_rom <= {16'd18428, 16'd27094};
                15'd6231 : data_rom <= {16'd18431, 16'd27092};
                15'd6232 : data_rom <= {16'd18434, 16'd27091};
                15'd6233 : data_rom <= {16'd18436, 16'd27089};
                15'd6234 : data_rom <= {16'd18439, 16'd27087};
                15'd6235 : data_rom <= {16'd18441, 16'd27085};
                15'd6236 : data_rom <= {16'd18444, 16'd27083};
                15'd6237 : data_rom <= {16'd18447, 16'd27082};
                15'd6238 : data_rom <= {16'd18449, 16'd27080};
                15'd6239 : data_rom <= {16'd18452, 16'd27078};
                15'd6240 : data_rom <= {16'd18454, 16'd27076};
                15'd6241 : data_rom <= {16'd18457, 16'd27075};
                15'd6242 : data_rom <= {16'd18460, 16'd27073};
                15'd6243 : data_rom <= {16'd18462, 16'd27071};
                15'd6244 : data_rom <= {16'd18465, 16'd27069};
                15'd6245 : data_rom <= {16'd18467, 16'd27068};
                15'd6246 : data_rom <= {16'd18470, 16'd27066};
                15'd6247 : data_rom <= {16'd18473, 16'd27064};
                15'd6248 : data_rom <= {16'd18475, 16'd27062};
                15'd6249 : data_rom <= {16'd18478, 16'd27060};
                15'd6250 : data_rom <= {16'd18480, 16'd27059};
                15'd6251 : data_rom <= {16'd18483, 16'd27057};
                15'd6252 : data_rom <= {16'd18486, 16'd27055};
                15'd6253 : data_rom <= {16'd18488, 16'd27053};
                15'd6254 : data_rom <= {16'd18491, 16'd27052};
                15'd6255 : data_rom <= {16'd18493, 16'd27050};
                15'd6256 : data_rom <= {16'd18496, 16'd27048};
                15'd6257 : data_rom <= {16'd18499, 16'd27046};
                15'd6258 : data_rom <= {16'd18501, 16'd27045};
                15'd6259 : data_rom <= {16'd18504, 16'd27043};
                15'd6260 : data_rom <= {16'd18506, 16'd27041};
                15'd6261 : data_rom <= {16'd18509, 16'd27039};
                15'd6262 : data_rom <= {16'd18511, 16'd27037};
                15'd6263 : data_rom <= {16'd18514, 16'd27036};
                15'd6264 : data_rom <= {16'd18517, 16'd27034};
                15'd6265 : data_rom <= {16'd18519, 16'd27032};
                15'd6266 : data_rom <= {16'd18522, 16'd27030};
                15'd6267 : data_rom <= {16'd18524, 16'd27029};
                15'd6268 : data_rom <= {16'd18527, 16'd27027};
                15'd6269 : data_rom <= {16'd18530, 16'd27025};
                15'd6270 : data_rom <= {16'd18532, 16'd27023};
                15'd6271 : data_rom <= {16'd18535, 16'd27021};
                15'd6272 : data_rom <= {16'd18537, 16'd27020};
                15'd6273 : data_rom <= {16'd18540, 16'd27018};
                15'd6274 : data_rom <= {16'd18543, 16'd27016};
                15'd6275 : data_rom <= {16'd18545, 16'd27014};
                15'd6276 : data_rom <= {16'd18548, 16'd27013};
                15'd6277 : data_rom <= {16'd18550, 16'd27011};
                15'd6278 : data_rom <= {16'd18553, 16'd27009};
                15'd6279 : data_rom <= {16'd18556, 16'd27007};
                15'd6280 : data_rom <= {16'd18558, 16'd27005};
                15'd6281 : data_rom <= {16'd18561, 16'd27004};
                15'd6282 : data_rom <= {16'd18563, 16'd27002};
                15'd6283 : data_rom <= {16'd18566, 16'd27000};
                15'd6284 : data_rom <= {16'd18568, 16'd26998};
                15'd6285 : data_rom <= {16'd18571, 16'd26997};
                15'd6286 : data_rom <= {16'd18574, 16'd26995};
                15'd6287 : data_rom <= {16'd18576, 16'd26993};
                15'd6288 : data_rom <= {16'd18579, 16'd26991};
                15'd6289 : data_rom <= {16'd18581, 16'd26989};
                15'd6290 : data_rom <= {16'd18584, 16'd26988};
                15'd6291 : data_rom <= {16'd18587, 16'd26986};
                15'd6292 : data_rom <= {16'd18589, 16'd26984};
                15'd6293 : data_rom <= {16'd18592, 16'd26982};
                15'd6294 : data_rom <= {16'd18594, 16'd26980};
                15'd6295 : data_rom <= {16'd18597, 16'd26979};
                15'd6296 : data_rom <= {16'd18600, 16'd26977};
                15'd6297 : data_rom <= {16'd18602, 16'd26975};
                15'd6298 : data_rom <= {16'd18605, 16'd26973};
                15'd6299 : data_rom <= {16'd18607, 16'd26972};
                15'd6300 : data_rom <= {16'd18610, 16'd26970};
                15'd6301 : data_rom <= {16'd18612, 16'd26968};
                15'd6302 : data_rom <= {16'd18615, 16'd26966};
                15'd6303 : data_rom <= {16'd18618, 16'd26964};
                15'd6304 : data_rom <= {16'd18620, 16'd26963};
                15'd6305 : data_rom <= {16'd18623, 16'd26961};
                15'd6306 : data_rom <= {16'd18625, 16'd26959};
                15'd6307 : data_rom <= {16'd18628, 16'd26957};
                15'd6308 : data_rom <= {16'd18631, 16'd26956};
                15'd6309 : data_rom <= {16'd18633, 16'd26954};
                15'd6310 : data_rom <= {16'd18636, 16'd26952};
                15'd6311 : data_rom <= {16'd18638, 16'd26950};
                15'd6312 : data_rom <= {16'd18641, 16'd26948};
                15'd6313 : data_rom <= {16'd18643, 16'd26947};
                15'd6314 : data_rom <= {16'd18646, 16'd26945};
                15'd6315 : data_rom <= {16'd18649, 16'd26943};
                15'd6316 : data_rom <= {16'd18651, 16'd26941};
                15'd6317 : data_rom <= {16'd18654, 16'd26939};
                15'd6318 : data_rom <= {16'd18656, 16'd26938};
                15'd6319 : data_rom <= {16'd18659, 16'd26936};
                15'd6320 : data_rom <= {16'd18662, 16'd26934};
                15'd6321 : data_rom <= {16'd18664, 16'd26932};
                15'd6322 : data_rom <= {16'd18667, 16'd26930};
                15'd6323 : data_rom <= {16'd18669, 16'd26929};
                15'd6324 : data_rom <= {16'd18672, 16'd26927};
                15'd6325 : data_rom <= {16'd18674, 16'd26925};
                15'd6326 : data_rom <= {16'd18677, 16'd26923};
                15'd6327 : data_rom <= {16'd18680, 16'd26922};
                15'd6328 : data_rom <= {16'd18682, 16'd26920};
                15'd6329 : data_rom <= {16'd18685, 16'd26918};
                15'd6330 : data_rom <= {16'd18687, 16'd26916};
                15'd6331 : data_rom <= {16'd18690, 16'd26914};
                15'd6332 : data_rom <= {16'd18693, 16'd26913};
                15'd6333 : data_rom <= {16'd18695, 16'd26911};
                15'd6334 : data_rom <= {16'd18698, 16'd26909};
                15'd6335 : data_rom <= {16'd18700, 16'd26907};
                15'd6336 : data_rom <= {16'd18703, 16'd26905};
                15'd6337 : data_rom <= {16'd18705, 16'd26904};
                15'd6338 : data_rom <= {16'd18708, 16'd26902};
                15'd6339 : data_rom <= {16'd18711, 16'd26900};
                15'd6340 : data_rom <= {16'd18713, 16'd26898};
                15'd6341 : data_rom <= {16'd18716, 16'd26896};
                15'd6342 : data_rom <= {16'd18718, 16'd26895};
                15'd6343 : data_rom <= {16'd18721, 16'd26893};
                15'd6344 : data_rom <= {16'd18723, 16'd26891};
                15'd6345 : data_rom <= {16'd18726, 16'd26889};
                15'd6346 : data_rom <= {16'd18729, 16'd26887};
                15'd6347 : data_rom <= {16'd18731, 16'd26886};
                15'd6348 : data_rom <= {16'd18734, 16'd26884};
                15'd6349 : data_rom <= {16'd18736, 16'd26882};
                15'd6350 : data_rom <= {16'd18739, 16'd26880};
                15'd6351 : data_rom <= {16'd18742, 16'd26878};
                15'd6352 : data_rom <= {16'd18744, 16'd26877};
                15'd6353 : data_rom <= {16'd18747, 16'd26875};
                15'd6354 : data_rom <= {16'd18749, 16'd26873};
                15'd6355 : data_rom <= {16'd18752, 16'd26871};
                15'd6356 : data_rom <= {16'd18754, 16'd26869};
                15'd6357 : data_rom <= {16'd18757, 16'd26868};
                15'd6358 : data_rom <= {16'd18760, 16'd26866};
                15'd6359 : data_rom <= {16'd18762, 16'd26864};
                15'd6360 : data_rom <= {16'd18765, 16'd26862};
                15'd6361 : data_rom <= {16'd18767, 16'd26860};
                15'd6362 : data_rom <= {16'd18770, 16'd26859};
                15'd6363 : data_rom <= {16'd18772, 16'd26857};
                15'd6364 : data_rom <= {16'd18775, 16'd26855};
                15'd6365 : data_rom <= {16'd18778, 16'd26853};
                15'd6366 : data_rom <= {16'd18780, 16'd26851};
                15'd6367 : data_rom <= {16'd18783, 16'd26850};
                15'd6368 : data_rom <= {16'd18785, 16'd26848};
                15'd6369 : data_rom <= {16'd18788, 16'd26846};
                15'd6370 : data_rom <= {16'd18790, 16'd26844};
                15'd6371 : data_rom <= {16'd18793, 16'd26842};
                15'd6372 : data_rom <= {16'd18796, 16'd26841};
                15'd6373 : data_rom <= {16'd18798, 16'd26839};
                15'd6374 : data_rom <= {16'd18801, 16'd26837};
                15'd6375 : data_rom <= {16'd18803, 16'd26835};
                15'd6376 : data_rom <= {16'd18806, 16'd26833};
                15'd6377 : data_rom <= {16'd18808, 16'd26832};
                15'd6378 : data_rom <= {16'd18811, 16'd26830};
                15'd6379 : data_rom <= {16'd18814, 16'd26828};
                15'd6380 : data_rom <= {16'd18816, 16'd26826};
                15'd6381 : data_rom <= {16'd18819, 16'd26824};
                15'd6382 : data_rom <= {16'd18821, 16'd26823};
                15'd6383 : data_rom <= {16'd18824, 16'd26821};
                15'd6384 : data_rom <= {16'd18826, 16'd26819};
                15'd6385 : data_rom <= {16'd18829, 16'd26817};
                15'd6386 : data_rom <= {16'd18832, 16'd26815};
                15'd6387 : data_rom <= {16'd18834, 16'd26814};
                15'd6388 : data_rom <= {16'd18837, 16'd26812};
                15'd6389 : data_rom <= {16'd18839, 16'd26810};
                15'd6390 : data_rom <= {16'd18842, 16'd26808};
                15'd6391 : data_rom <= {16'd18844, 16'd26806};
                15'd6392 : data_rom <= {16'd18847, 16'd26805};
                15'd6393 : data_rom <= {16'd18850, 16'd26803};
                15'd6394 : data_rom <= {16'd18852, 16'd26801};
                15'd6395 : data_rom <= {16'd18855, 16'd26799};
                15'd6396 : data_rom <= {16'd18857, 16'd26797};
                15'd6397 : data_rom <= {16'd18860, 16'd26796};
                15'd6398 : data_rom <= {16'd18862, 16'd26794};
                15'd6399 : data_rom <= {16'd18865, 16'd26792};
                15'd6400 : data_rom <= {16'd18868, 16'd26790};
                15'd6401 : data_rom <= {16'd18870, 16'd26788};
                15'd6402 : data_rom <= {16'd18873, 16'd26787};
                15'd6403 : data_rom <= {16'd18875, 16'd26785};
                15'd6404 : data_rom <= {16'd18878, 16'd26783};
                15'd6405 : data_rom <= {16'd18880, 16'd26781};
                15'd6406 : data_rom <= {16'd18883, 16'd26779};
                15'd6407 : data_rom <= {16'd18886, 16'd26777};
                15'd6408 : data_rom <= {16'd18888, 16'd26776};
                15'd6409 : data_rom <= {16'd18891, 16'd26774};
                15'd6410 : data_rom <= {16'd18893, 16'd26772};
                15'd6411 : data_rom <= {16'd18896, 16'd26770};
                15'd6412 : data_rom <= {16'd18898, 16'd26768};
                15'd6413 : data_rom <= {16'd18901, 16'd26767};
                15'd6414 : data_rom <= {16'd18904, 16'd26765};
                15'd6415 : data_rom <= {16'd18906, 16'd26763};
                15'd6416 : data_rom <= {16'd18909, 16'd26761};
                15'd6417 : data_rom <= {16'd18911, 16'd26759};
                15'd6418 : data_rom <= {16'd18914, 16'd26758};
                15'd6419 : data_rom <= {16'd18916, 16'd26756};
                15'd6420 : data_rom <= {16'd18919, 16'd26754};
                15'd6421 : data_rom <= {16'd18921, 16'd26752};
                15'd6422 : data_rom <= {16'd18924, 16'd26750};
                15'd6423 : data_rom <= {16'd18927, 16'd26748};
                15'd6424 : data_rom <= {16'd18929, 16'd26747};
                15'd6425 : data_rom <= {16'd18932, 16'd26745};
                15'd6426 : data_rom <= {16'd18934, 16'd26743};
                15'd6427 : data_rom <= {16'd18937, 16'd26741};
                15'd6428 : data_rom <= {16'd18939, 16'd26739};
                15'd6429 : data_rom <= {16'd18942, 16'd26738};
                15'd6430 : data_rom <= {16'd18945, 16'd26736};
                15'd6431 : data_rom <= {16'd18947, 16'd26734};
                15'd6432 : data_rom <= {16'd18950, 16'd26732};
                15'd6433 : data_rom <= {16'd18952, 16'd26730};
                15'd6434 : data_rom <= {16'd18955, 16'd26728};
                15'd6435 : data_rom <= {16'd18957, 16'd26727};
                15'd6436 : data_rom <= {16'd18960, 16'd26725};
                15'd6437 : data_rom <= {16'd18962, 16'd26723};
                15'd6438 : data_rom <= {16'd18965, 16'd26721};
                15'd6439 : data_rom <= {16'd18968, 16'd26719};
                15'd6440 : data_rom <= {16'd18970, 16'd26718};
                15'd6441 : data_rom <= {16'd18973, 16'd26716};
                15'd6442 : data_rom <= {16'd18975, 16'd26714};
                15'd6443 : data_rom <= {16'd18978, 16'd26712};
                15'd6444 : data_rom <= {16'd18980, 16'd26710};
                15'd6445 : data_rom <= {16'd18983, 16'd26708};
                15'd6446 : data_rom <= {16'd18986, 16'd26707};
                15'd6447 : data_rom <= {16'd18988, 16'd26705};
                15'd6448 : data_rom <= {16'd18991, 16'd26703};
                15'd6449 : data_rom <= {16'd18993, 16'd26701};
                15'd6450 : data_rom <= {16'd18996, 16'd26699};
                15'd6451 : data_rom <= {16'd18998, 16'd26698};
                15'd6452 : data_rom <= {16'd19001, 16'd26696};
                15'd6453 : data_rom <= {16'd19003, 16'd26694};
                15'd6454 : data_rom <= {16'd19006, 16'd26692};
                15'd6455 : data_rom <= {16'd19009, 16'd26690};
                15'd6456 : data_rom <= {16'd19011, 16'd26688};
                15'd6457 : data_rom <= {16'd19014, 16'd26687};
                15'd6458 : data_rom <= {16'd19016, 16'd26685};
                15'd6459 : data_rom <= {16'd19019, 16'd26683};
                15'd6460 : data_rom <= {16'd19021, 16'd26681};
                15'd6461 : data_rom <= {16'd19024, 16'd26679};
                15'd6462 : data_rom <= {16'd19026, 16'd26678};
                15'd6463 : data_rom <= {16'd19029, 16'd26676};
                15'd6464 : data_rom <= {16'd19032, 16'd26674};
                15'd6465 : data_rom <= {16'd19034, 16'd26672};
                15'd6466 : data_rom <= {16'd19037, 16'd26670};
                15'd6467 : data_rom <= {16'd19039, 16'd26668};
                15'd6468 : data_rom <= {16'd19042, 16'd26667};
                15'd6469 : data_rom <= {16'd19044, 16'd26665};
                15'd6470 : data_rom <= {16'd19047, 16'd26663};
                15'd6471 : data_rom <= {16'd19049, 16'd26661};
                15'd6472 : data_rom <= {16'd19052, 16'd26659};
                15'd6473 : data_rom <= {16'd19055, 16'd26657};
                15'd6474 : data_rom <= {16'd19057, 16'd26656};
                15'd6475 : data_rom <= {16'd19060, 16'd26654};
                15'd6476 : data_rom <= {16'd19062, 16'd26652};
                15'd6477 : data_rom <= {16'd19065, 16'd26650};
                15'd6478 : data_rom <= {16'd19067, 16'd26648};
                15'd6479 : data_rom <= {16'd19070, 16'd26646};
                15'd6480 : data_rom <= {16'd19072, 16'd26645};
                15'd6481 : data_rom <= {16'd19075, 16'd26643};
                15'd6482 : data_rom <= {16'd19078, 16'd26641};
                15'd6483 : data_rom <= {16'd19080, 16'd26639};
                15'd6484 : data_rom <= {16'd19083, 16'd26637};
                15'd6485 : data_rom <= {16'd19085, 16'd26635};
                15'd6486 : data_rom <= {16'd19088, 16'd26634};
                15'd6487 : data_rom <= {16'd19090, 16'd26632};
                15'd6488 : data_rom <= {16'd19093, 16'd26630};
                15'd6489 : data_rom <= {16'd19095, 16'd26628};
                15'd6490 : data_rom <= {16'd19098, 16'd26626};
                15'd6491 : data_rom <= {16'd19101, 16'd26624};
                15'd6492 : data_rom <= {16'd19103, 16'd26623};
                15'd6493 : data_rom <= {16'd19106, 16'd26621};
                15'd6494 : data_rom <= {16'd19108, 16'd26619};
                15'd6495 : data_rom <= {16'd19111, 16'd26617};
                15'd6496 : data_rom <= {16'd19113, 16'd26615};
                15'd6497 : data_rom <= {16'd19116, 16'd26614};
                15'd6498 : data_rom <= {16'd19118, 16'd26612};
                15'd6499 : data_rom <= {16'd19121, 16'd26610};
                15'd6500 : data_rom <= {16'd19124, 16'd26608};
                15'd6501 : data_rom <= {16'd19126, 16'd26606};
                15'd6502 : data_rom <= {16'd19129, 16'd26604};
                15'd6503 : data_rom <= {16'd19131, 16'd26603};
                15'd6504 : data_rom <= {16'd19134, 16'd26601};
                15'd6505 : data_rom <= {16'd19136, 16'd26599};
                15'd6506 : data_rom <= {16'd19139, 16'd26597};
                15'd6507 : data_rom <= {16'd19141, 16'd26595};
                15'd6508 : data_rom <= {16'd19144, 16'd26593};
                15'd6509 : data_rom <= {16'd19147, 16'd26591};
                15'd6510 : data_rom <= {16'd19149, 16'd26590};
                15'd6511 : data_rom <= {16'd19152, 16'd26588};
                15'd6512 : data_rom <= {16'd19154, 16'd26586};
                15'd6513 : data_rom <= {16'd19157, 16'd26584};
                15'd6514 : data_rom <= {16'd19159, 16'd26582};
                15'd6515 : data_rom <= {16'd19162, 16'd26580};
                15'd6516 : data_rom <= {16'd19164, 16'd26579};
                15'd6517 : data_rom <= {16'd19167, 16'd26577};
                15'd6518 : data_rom <= {16'd19169, 16'd26575};
                15'd6519 : data_rom <= {16'd19172, 16'd26573};
                15'd6520 : data_rom <= {16'd19175, 16'd26571};
                15'd6521 : data_rom <= {16'd19177, 16'd26569};
                15'd6522 : data_rom <= {16'd19180, 16'd26568};
                15'd6523 : data_rom <= {16'd19182, 16'd26566};
                15'd6524 : data_rom <= {16'd19185, 16'd26564};
                15'd6525 : data_rom <= {16'd19187, 16'd26562};
                15'd6526 : data_rom <= {16'd19190, 16'd26560};
                15'd6527 : data_rom <= {16'd19192, 16'd26558};
                15'd6528 : data_rom <= {16'd19195, 16'd26557};
                15'd6529 : data_rom <= {16'd19197, 16'd26555};
                15'd6530 : data_rom <= {16'd19200, 16'd26553};
                15'd6531 : data_rom <= {16'd19203, 16'd26551};
                15'd6532 : data_rom <= {16'd19205, 16'd26549};
                15'd6533 : data_rom <= {16'd19208, 16'd26547};
                15'd6534 : data_rom <= {16'd19210, 16'd26546};
                15'd6535 : data_rom <= {16'd19213, 16'd26544};
                15'd6536 : data_rom <= {16'd19215, 16'd26542};
                15'd6537 : data_rom <= {16'd19218, 16'd26540};
                15'd6538 : data_rom <= {16'd19220, 16'd26538};
                15'd6539 : data_rom <= {16'd19223, 16'd26536};
                15'd6540 : data_rom <= {16'd19225, 16'd26534};
                15'd6541 : data_rom <= {16'd19228, 16'd26533};
                15'd6542 : data_rom <= {16'd19231, 16'd26531};
                15'd6543 : data_rom <= {16'd19233, 16'd26529};
                15'd6544 : data_rom <= {16'd19236, 16'd26527};
                15'd6545 : data_rom <= {16'd19238, 16'd26525};
                15'd6546 : data_rom <= {16'd19241, 16'd26523};
                15'd6547 : data_rom <= {16'd19243, 16'd26522};
                15'd6548 : data_rom <= {16'd19246, 16'd26520};
                15'd6549 : data_rom <= {16'd19248, 16'd26518};
                15'd6550 : data_rom <= {16'd19251, 16'd26516};
                15'd6551 : data_rom <= {16'd19253, 16'd26514};
                15'd6552 : data_rom <= {16'd19256, 16'd26512};
                15'd6553 : data_rom <= {16'd19259, 16'd26510};
                15'd6554 : data_rom <= {16'd19261, 16'd26509};
                15'd6555 : data_rom <= {16'd19264, 16'd26507};
                15'd6556 : data_rom <= {16'd19266, 16'd26505};
                15'd6557 : data_rom <= {16'd19269, 16'd26503};
                15'd6558 : data_rom <= {16'd19271, 16'd26501};
                15'd6559 : data_rom <= {16'd19274, 16'd26499};
                15'd6560 : data_rom <= {16'd19276, 16'd26498};
                15'd6561 : data_rom <= {16'd19279, 16'd26496};
                15'd6562 : data_rom <= {16'd19281, 16'd26494};
                15'd6563 : data_rom <= {16'd19284, 16'd26492};
                15'd6564 : data_rom <= {16'd19286, 16'd26490};
                15'd6565 : data_rom <= {16'd19289, 16'd26488};
                15'd6566 : data_rom <= {16'd19292, 16'd26486};
                15'd6567 : data_rom <= {16'd19294, 16'd26485};
                15'd6568 : data_rom <= {16'd19297, 16'd26483};
                15'd6569 : data_rom <= {16'd19299, 16'd26481};
                15'd6570 : data_rom <= {16'd19302, 16'd26479};
                15'd6571 : data_rom <= {16'd19304, 16'd26477};
                15'd6572 : data_rom <= {16'd19307, 16'd26475};
                15'd6573 : data_rom <= {16'd19309, 16'd26474};
                15'd6574 : data_rom <= {16'd19312, 16'd26472};
                15'd6575 : data_rom <= {16'd19314, 16'd26470};
                15'd6576 : data_rom <= {16'd19317, 16'd26468};
                15'd6577 : data_rom <= {16'd19319, 16'd26466};
                15'd6578 : data_rom <= {16'd19322, 16'd26464};
                15'd6579 : data_rom <= {16'd19325, 16'd26462};
                15'd6580 : data_rom <= {16'd19327, 16'd26461};
                15'd6581 : data_rom <= {16'd19330, 16'd26459};
                15'd6582 : data_rom <= {16'd19332, 16'd26457};
                15'd6583 : data_rom <= {16'd19335, 16'd26455};
                15'd6584 : data_rom <= {16'd19337, 16'd26453};
                15'd6585 : data_rom <= {16'd19340, 16'd26451};
                15'd6586 : data_rom <= {16'd19342, 16'd26449};
                15'd6587 : data_rom <= {16'd19345, 16'd26448};
                15'd6588 : data_rom <= {16'd19347, 16'd26446};
                15'd6589 : data_rom <= {16'd19350, 16'd26444};
                15'd6590 : data_rom <= {16'd19352, 16'd26442};
                15'd6591 : data_rom <= {16'd19355, 16'd26440};
                15'd6592 : data_rom <= {16'd19357, 16'd26438};
                15'd6593 : data_rom <= {16'd19360, 16'd26436};
                15'd6594 : data_rom <= {16'd19363, 16'd26435};
                15'd6595 : data_rom <= {16'd19365, 16'd26433};
                15'd6596 : data_rom <= {16'd19368, 16'd26431};
                15'd6597 : data_rom <= {16'd19370, 16'd26429};
                15'd6598 : data_rom <= {16'd19373, 16'd26427};
                15'd6599 : data_rom <= {16'd19375, 16'd26425};
                15'd6600 : data_rom <= {16'd19378, 16'd26423};
                15'd6601 : data_rom <= {16'd19380, 16'd26422};
                15'd6602 : data_rom <= {16'd19383, 16'd26420};
                15'd6603 : data_rom <= {16'd19385, 16'd26418};
                15'd6604 : data_rom <= {16'd19388, 16'd26416};
                15'd6605 : data_rom <= {16'd19390, 16'd26414};
                15'd6606 : data_rom <= {16'd19393, 16'd26412};
                15'd6607 : data_rom <= {16'd19395, 16'd26410};
                15'd6608 : data_rom <= {16'd19398, 16'd26409};
                15'd6609 : data_rom <= {16'd19401, 16'd26407};
                15'd6610 : data_rom <= {16'd19403, 16'd26405};
                15'd6611 : data_rom <= {16'd19406, 16'd26403};
                15'd6612 : data_rom <= {16'd19408, 16'd26401};
                15'd6613 : data_rom <= {16'd19411, 16'd26399};
                15'd6614 : data_rom <= {16'd19413, 16'd26397};
                15'd6615 : data_rom <= {16'd19416, 16'd26396};
                15'd6616 : data_rom <= {16'd19418, 16'd26394};
                15'd6617 : data_rom <= {16'd19421, 16'd26392};
                15'd6618 : data_rom <= {16'd19423, 16'd26390};
                15'd6619 : data_rom <= {16'd19426, 16'd26388};
                15'd6620 : data_rom <= {16'd19428, 16'd26386};
                15'd6621 : data_rom <= {16'd19431, 16'd26384};
                15'd6622 : data_rom <= {16'd19433, 16'd26383};
                15'd6623 : data_rom <= {16'd19436, 16'd26381};
                15'd6624 : data_rom <= {16'd19439, 16'd26379};
                15'd6625 : data_rom <= {16'd19441, 16'd26377};
                15'd6626 : data_rom <= {16'd19444, 16'd26375};
                15'd6627 : data_rom <= {16'd19446, 16'd26373};
                15'd6628 : data_rom <= {16'd19449, 16'd26371};
                15'd6629 : data_rom <= {16'd19451, 16'd26369};
                15'd6630 : data_rom <= {16'd19454, 16'd26368};
                15'd6631 : data_rom <= {16'd19456, 16'd26366};
                15'd6632 : data_rom <= {16'd19459, 16'd26364};
                15'd6633 : data_rom <= {16'd19461, 16'd26362};
                15'd6634 : data_rom <= {16'd19464, 16'd26360};
                15'd6635 : data_rom <= {16'd19466, 16'd26358};
                15'd6636 : data_rom <= {16'd19469, 16'd26356};
                15'd6637 : data_rom <= {16'd19471, 16'd26355};
                15'd6638 : data_rom <= {16'd19474, 16'd26353};
                15'd6639 : data_rom <= {16'd19476, 16'd26351};
                15'd6640 : data_rom <= {16'd19479, 16'd26349};
                15'd6641 : data_rom <= {16'd19481, 16'd26347};
                15'd6642 : data_rom <= {16'd19484, 16'd26345};
                15'd6643 : data_rom <= {16'd19487, 16'd26343};
                15'd6644 : data_rom <= {16'd19489, 16'd26341};
                15'd6645 : data_rom <= {16'd19492, 16'd26340};
                15'd6646 : data_rom <= {16'd19494, 16'd26338};
                15'd6647 : data_rom <= {16'd19497, 16'd26336};
                15'd6648 : data_rom <= {16'd19499, 16'd26334};
                15'd6649 : data_rom <= {16'd19502, 16'd26332};
                15'd6650 : data_rom <= {16'd19504, 16'd26330};
                15'd6651 : data_rom <= {16'd19507, 16'd26328};
                15'd6652 : data_rom <= {16'd19509, 16'd26327};
                15'd6653 : data_rom <= {16'd19512, 16'd26325};
                15'd6654 : data_rom <= {16'd19514, 16'd26323};
                15'd6655 : data_rom <= {16'd19517, 16'd26321};
                15'd6656 : data_rom <= {16'd19519, 16'd26319};
                15'd6657 : data_rom <= {16'd19522, 16'd26317};
                15'd6658 : data_rom <= {16'd19524, 16'd26315};
                15'd6659 : data_rom <= {16'd19527, 16'd26313};
                15'd6660 : data_rom <= {16'd19529, 16'd26312};
                15'd6661 : data_rom <= {16'd19532, 16'd26310};
                15'd6662 : data_rom <= {16'd19534, 16'd26308};
                15'd6663 : data_rom <= {16'd19537, 16'd26306};
                15'd6664 : data_rom <= {16'd19540, 16'd26304};
                15'd6665 : data_rom <= {16'd19542, 16'd26302};
                15'd6666 : data_rom <= {16'd19545, 16'd26300};
                15'd6667 : data_rom <= {16'd19547, 16'd26298};
                15'd6668 : data_rom <= {16'd19550, 16'd26297};
                15'd6669 : data_rom <= {16'd19552, 16'd26295};
                15'd6670 : data_rom <= {16'd19555, 16'd26293};
                15'd6671 : data_rom <= {16'd19557, 16'd26291};
                15'd6672 : data_rom <= {16'd19560, 16'd26289};
                15'd6673 : data_rom <= {16'd19562, 16'd26287};
                15'd6674 : data_rom <= {16'd19565, 16'd26285};
                15'd6675 : data_rom <= {16'd19567, 16'd26283};
                15'd6676 : data_rom <= {16'd19570, 16'd26282};
                15'd6677 : data_rom <= {16'd19572, 16'd26280};
                15'd6678 : data_rom <= {16'd19575, 16'd26278};
                15'd6679 : data_rom <= {16'd19577, 16'd26276};
                15'd6680 : data_rom <= {16'd19580, 16'd26274};
                15'd6681 : data_rom <= {16'd19582, 16'd26272};
                15'd6682 : data_rom <= {16'd19585, 16'd26270};
                15'd6683 : data_rom <= {16'd19587, 16'd26268};
                15'd6684 : data_rom <= {16'd19590, 16'd26267};
                15'd6685 : data_rom <= {16'd19592, 16'd26265};
                15'd6686 : data_rom <= {16'd19595, 16'd26263};
                15'd6687 : data_rom <= {16'd19597, 16'd26261};
                15'd6688 : data_rom <= {16'd19600, 16'd26259};
                15'd6689 : data_rom <= {16'd19603, 16'd26257};
                15'd6690 : data_rom <= {16'd19605, 16'd26255};
                15'd6691 : data_rom <= {16'd19608, 16'd26253};
                15'd6692 : data_rom <= {16'd19610, 16'd26251};
                15'd6693 : data_rom <= {16'd19613, 16'd26250};
                15'd6694 : data_rom <= {16'd19615, 16'd26248};
                15'd6695 : data_rom <= {16'd19618, 16'd26246};
                15'd6696 : data_rom <= {16'd19620, 16'd26244};
                15'd6697 : data_rom <= {16'd19623, 16'd26242};
                15'd6698 : data_rom <= {16'd19625, 16'd26240};
                15'd6699 : data_rom <= {16'd19628, 16'd26238};
                15'd6700 : data_rom <= {16'd19630, 16'd26236};
                15'd6701 : data_rom <= {16'd19633, 16'd26235};
                15'd6702 : data_rom <= {16'd19635, 16'd26233};
                15'd6703 : data_rom <= {16'd19638, 16'd26231};
                15'd6704 : data_rom <= {16'd19640, 16'd26229};
                15'd6705 : data_rom <= {16'd19643, 16'd26227};
                15'd6706 : data_rom <= {16'd19645, 16'd26225};
                15'd6707 : data_rom <= {16'd19648, 16'd26223};
                15'd6708 : data_rom <= {16'd19650, 16'd26221};
                15'd6709 : data_rom <= {16'd19653, 16'd26219};
                15'd6710 : data_rom <= {16'd19655, 16'd26218};
                15'd6711 : data_rom <= {16'd19658, 16'd26216};
                15'd6712 : data_rom <= {16'd19660, 16'd26214};
                15'd6713 : data_rom <= {16'd19663, 16'd26212};
                15'd6714 : data_rom <= {16'd19665, 16'd26210};
                15'd6715 : data_rom <= {16'd19668, 16'd26208};
                15'd6716 : data_rom <= {16'd19670, 16'd26206};
                15'd6717 : data_rom <= {16'd19673, 16'd26204};
                15'd6718 : data_rom <= {16'd19675, 16'd26203};
                15'd6719 : data_rom <= {16'd19678, 16'd26201};
                15'd6720 : data_rom <= {16'd19680, 16'd26199};
                15'd6721 : data_rom <= {16'd19683, 16'd26197};
                15'd6722 : data_rom <= {16'd19686, 16'd26195};
                15'd6723 : data_rom <= {16'd19688, 16'd26193};
                15'd6724 : data_rom <= {16'd19691, 16'd26191};
                15'd6725 : data_rom <= {16'd19693, 16'd26189};
                15'd6726 : data_rom <= {16'd19696, 16'd26187};
                15'd6727 : data_rom <= {16'd19698, 16'd26186};
                15'd6728 : data_rom <= {16'd19701, 16'd26184};
                15'd6729 : data_rom <= {16'd19703, 16'd26182};
                15'd6730 : data_rom <= {16'd19706, 16'd26180};
                15'd6731 : data_rom <= {16'd19708, 16'd26178};
                15'd6732 : data_rom <= {16'd19711, 16'd26176};
                15'd6733 : data_rom <= {16'd19713, 16'd26174};
                15'd6734 : data_rom <= {16'd19716, 16'd26172};
                15'd6735 : data_rom <= {16'd19718, 16'd26170};
                15'd6736 : data_rom <= {16'd19721, 16'd26169};
                15'd6737 : data_rom <= {16'd19723, 16'd26167};
                15'd6738 : data_rom <= {16'd19726, 16'd26165};
                15'd6739 : data_rom <= {16'd19728, 16'd26163};
                15'd6740 : data_rom <= {16'd19731, 16'd26161};
                15'd6741 : data_rom <= {16'd19733, 16'd26159};
                15'd6742 : data_rom <= {16'd19736, 16'd26157};
                15'd6743 : data_rom <= {16'd19738, 16'd26155};
                15'd6744 : data_rom <= {16'd19741, 16'd26153};
                15'd6745 : data_rom <= {16'd19743, 16'd26152};
                15'd6746 : data_rom <= {16'd19746, 16'd26150};
                15'd6747 : data_rom <= {16'd19748, 16'd26148};
                15'd6748 : data_rom <= {16'd19751, 16'd26146};
                15'd6749 : data_rom <= {16'd19753, 16'd26144};
                15'd6750 : data_rom <= {16'd19756, 16'd26142};
                15'd6751 : data_rom <= {16'd19758, 16'd26140};
                15'd6752 : data_rom <= {16'd19761, 16'd26138};
                15'd6753 : data_rom <= {16'd19763, 16'd26136};
                15'd6754 : data_rom <= {16'd19766, 16'd26134};
                15'd6755 : data_rom <= {16'd19768, 16'd26133};
                15'd6756 : data_rom <= {16'd19771, 16'd26131};
                15'd6757 : data_rom <= {16'd19773, 16'd26129};
                15'd6758 : data_rom <= {16'd19776, 16'd26127};
                15'd6759 : data_rom <= {16'd19778, 16'd26125};
                15'd6760 : data_rom <= {16'd19781, 16'd26123};
                15'd6761 : data_rom <= {16'd19783, 16'd26121};
                15'd6762 : data_rom <= {16'd19786, 16'd26119};
                15'd6763 : data_rom <= {16'd19788, 16'd26117};
                15'd6764 : data_rom <= {16'd19791, 16'd26115};
                15'd6765 : data_rom <= {16'd19793, 16'd26114};
                15'd6766 : data_rom <= {16'd19796, 16'd26112};
                15'd6767 : data_rom <= {16'd19798, 16'd26110};
                15'd6768 : data_rom <= {16'd19801, 16'd26108};
                15'd6769 : data_rom <= {16'd19803, 16'd26106};
                15'd6770 : data_rom <= {16'd19806, 16'd26104};
                15'd6771 : data_rom <= {16'd19808, 16'd26102};
                15'd6772 : data_rom <= {16'd19811, 16'd26100};
                15'd6773 : data_rom <= {16'd19813, 16'd26098};
                15'd6774 : data_rom <= {16'd19816, 16'd26097};
                15'd6775 : data_rom <= {16'd19818, 16'd26095};
                15'd6776 : data_rom <= {16'd19821, 16'd26093};
                15'd6777 : data_rom <= {16'd19823, 16'd26091};
                15'd6778 : data_rom <= {16'd19826, 16'd26089};
                15'd6779 : data_rom <= {16'd19828, 16'd26087};
                15'd6780 : data_rom <= {16'd19831, 16'd26085};
                15'd6781 : data_rom <= {16'd19833, 16'd26083};
                15'd6782 : data_rom <= {16'd19836, 16'd26081};
                15'd6783 : data_rom <= {16'd19838, 16'd26079};
                15'd6784 : data_rom <= {16'd19841, 16'd26077};
                15'd6785 : data_rom <= {16'd19843, 16'd26076};
                15'd6786 : data_rom <= {16'd19846, 16'd26074};
                15'd6787 : data_rom <= {16'd19848, 16'd26072};
                15'd6788 : data_rom <= {16'd19851, 16'd26070};
                15'd6789 : data_rom <= {16'd19853, 16'd26068};
                15'd6790 : data_rom <= {16'd19856, 16'd26066};
                15'd6791 : data_rom <= {16'd19858, 16'd26064};
                15'd6792 : data_rom <= {16'd19861, 16'd26062};
                15'd6793 : data_rom <= {16'd19863, 16'd26060};
                15'd6794 : data_rom <= {16'd19866, 16'd26058};
                15'd6795 : data_rom <= {16'd19868, 16'd26057};
                15'd6796 : data_rom <= {16'd19871, 16'd26055};
                15'd6797 : data_rom <= {16'd19873, 16'd26053};
                15'd6798 : data_rom <= {16'd19876, 16'd26051};
                15'd6799 : data_rom <= {16'd19878, 16'd26049};
                15'd6800 : data_rom <= {16'd19881, 16'd26047};
                15'd6801 : data_rom <= {16'd19883, 16'd26045};
                15'd6802 : data_rom <= {16'd19886, 16'd26043};
                15'd6803 : data_rom <= {16'd19888, 16'd26041};
                15'd6804 : data_rom <= {16'd19891, 16'd26039};
                15'd6805 : data_rom <= {16'd19893, 16'd26037};
                15'd6806 : data_rom <= {16'd19896, 16'd26036};
                15'd6807 : data_rom <= {16'd19898, 16'd26034};
                15'd6808 : data_rom <= {16'd19901, 16'd26032};
                15'd6809 : data_rom <= {16'd19903, 16'd26030};
                15'd6810 : data_rom <= {16'd19906, 16'd26028};
                15'd6811 : data_rom <= {16'd19908, 16'd26026};
                15'd6812 : data_rom <= {16'd19911, 16'd26024};
                15'd6813 : data_rom <= {16'd19913, 16'd26022};
                15'd6814 : data_rom <= {16'd19916, 16'd26020};
                15'd6815 : data_rom <= {16'd19918, 16'd26018};
                15'd6816 : data_rom <= {16'd19921, 16'd26017};
                15'd6817 : data_rom <= {16'd19923, 16'd26015};
                15'd6818 : data_rom <= {16'd19926, 16'd26013};
                15'd6819 : data_rom <= {16'd19928, 16'd26011};
                15'd6820 : data_rom <= {16'd19931, 16'd26009};
                15'd6821 : data_rom <= {16'd19933, 16'd26007};
                15'd6822 : data_rom <= {16'd19936, 16'd26005};
                15'd6823 : data_rom <= {16'd19938, 16'd26003};
                15'd6824 : data_rom <= {16'd19941, 16'd26001};
                15'd6825 : data_rom <= {16'd19943, 16'd25999};
                15'd6826 : data_rom <= {16'd19946, 16'd25997};
                15'd6827 : data_rom <= {16'd19948, 16'd25995};
                15'd6828 : data_rom <= {16'd19951, 16'd25994};
                15'd6829 : data_rom <= {16'd19953, 16'd25992};
                15'd6830 : data_rom <= {16'd19956, 16'd25990};
                15'd6831 : data_rom <= {16'd19958, 16'd25988};
                15'd6832 : data_rom <= {16'd19961, 16'd25986};
                15'd6833 : data_rom <= {16'd19963, 16'd25984};
                15'd6834 : data_rom <= {16'd19966, 16'd25982};
                15'd6835 : data_rom <= {16'd19968, 16'd25980};
                15'd6836 : data_rom <= {16'd19971, 16'd25978};
                15'd6837 : data_rom <= {16'd19973, 16'd25976};
                15'd6838 : data_rom <= {16'd19976, 16'd25974};
                15'd6839 : data_rom <= {16'd19978, 16'd25973};
                15'd6840 : data_rom <= {16'd19981, 16'd25971};
                15'd6841 : data_rom <= {16'd19983, 16'd25969};
                15'd6842 : data_rom <= {16'd19986, 16'd25967};
                15'd6843 : data_rom <= {16'd19988, 16'd25965};
                15'd6844 : data_rom <= {16'd19991, 16'd25963};
                15'd6845 : data_rom <= {16'd19993, 16'd25961};
                15'd6846 : data_rom <= {16'd19996, 16'd25959};
                15'd6847 : data_rom <= {16'd19998, 16'd25957};
                15'd6848 : data_rom <= {16'd20001, 16'd25955};
                15'd6849 : data_rom <= {16'd20003, 16'd25953};
                15'd6850 : data_rom <= {16'd20005, 16'd25951};
                15'd6851 : data_rom <= {16'd20008, 16'd25950};
                15'd6852 : data_rom <= {16'd20010, 16'd25948};
                15'd6853 : data_rom <= {16'd20013, 16'd25946};
                15'd6854 : data_rom <= {16'd20015, 16'd25944};
                15'd6855 : data_rom <= {16'd20018, 16'd25942};
                15'd6856 : data_rom <= {16'd20020, 16'd25940};
                15'd6857 : data_rom <= {16'd20023, 16'd25938};
                15'd6858 : data_rom <= {16'd20025, 16'd25936};
                15'd6859 : data_rom <= {16'd20028, 16'd25934};
                15'd6860 : data_rom <= {16'd20030, 16'd25932};
                15'd6861 : data_rom <= {16'd20033, 16'd25930};
                15'd6862 : data_rom <= {16'd20035, 16'd25928};
                15'd6863 : data_rom <= {16'd20038, 16'd25926};
                15'd6864 : data_rom <= {16'd20040, 16'd25925};
                15'd6865 : data_rom <= {16'd20043, 16'd25923};
                15'd6866 : data_rom <= {16'd20045, 16'd25921};
                15'd6867 : data_rom <= {16'd20048, 16'd25919};
                15'd6868 : data_rom <= {16'd20050, 16'd25917};
                15'd6869 : data_rom <= {16'd20053, 16'd25915};
                15'd6870 : data_rom <= {16'd20055, 16'd25913};
                15'd6871 : data_rom <= {16'd20058, 16'd25911};
                15'd6872 : data_rom <= {16'd20060, 16'd25909};
                15'd6873 : data_rom <= {16'd20063, 16'd25907};
                15'd6874 : data_rom <= {16'd20065, 16'd25905};
                15'd6875 : data_rom <= {16'd20068, 16'd25903};
                15'd6876 : data_rom <= {16'd20070, 16'd25901};
                15'd6877 : data_rom <= {16'd20073, 16'd25900};
                15'd6878 : data_rom <= {16'd20075, 16'd25898};
                15'd6879 : data_rom <= {16'd20078, 16'd25896};
                15'd6880 : data_rom <= {16'd20080, 16'd25894};
                15'd6881 : data_rom <= {16'd20083, 16'd25892};
                15'd6882 : data_rom <= {16'd20085, 16'd25890};
                15'd6883 : data_rom <= {16'd20087, 16'd25888};
                15'd6884 : data_rom <= {16'd20090, 16'd25886};
                15'd6885 : data_rom <= {16'd20092, 16'd25884};
                15'd6886 : data_rom <= {16'd20095, 16'd25882};
                15'd6887 : data_rom <= {16'd20097, 16'd25880};
                15'd6888 : data_rom <= {16'd20100, 16'd25878};
                15'd6889 : data_rom <= {16'd20102, 16'd25876};
                15'd6890 : data_rom <= {16'd20105, 16'd25875};
                15'd6891 : data_rom <= {16'd20107, 16'd25873};
                15'd6892 : data_rom <= {16'd20110, 16'd25871};
                15'd6893 : data_rom <= {16'd20112, 16'd25869};
                15'd6894 : data_rom <= {16'd20115, 16'd25867};
                15'd6895 : data_rom <= {16'd20117, 16'd25865};
                15'd6896 : data_rom <= {16'd20120, 16'd25863};
                15'd6897 : data_rom <= {16'd20122, 16'd25861};
                15'd6898 : data_rom <= {16'd20125, 16'd25859};
                15'd6899 : data_rom <= {16'd20127, 16'd25857};
                15'd6900 : data_rom <= {16'd20130, 16'd25855};
                15'd6901 : data_rom <= {16'd20132, 16'd25853};
                15'd6902 : data_rom <= {16'd20135, 16'd25851};
                15'd6903 : data_rom <= {16'd20137, 16'd25849};
                15'd6904 : data_rom <= {16'd20140, 16'd25848};
                15'd6905 : data_rom <= {16'd20142, 16'd25846};
                15'd6906 : data_rom <= {16'd20145, 16'd25844};
                15'd6907 : data_rom <= {16'd20147, 16'd25842};
                15'd6908 : data_rom <= {16'd20149, 16'd25840};
                15'd6909 : data_rom <= {16'd20152, 16'd25838};
                15'd6910 : data_rom <= {16'd20154, 16'd25836};
                15'd6911 : data_rom <= {16'd20157, 16'd25834};
                15'd6912 : data_rom <= {16'd20159, 16'd25832};
                15'd6913 : data_rom <= {16'd20162, 16'd25830};
                15'd6914 : data_rom <= {16'd20164, 16'd25828};
                15'd6915 : data_rom <= {16'd20167, 16'd25826};
                15'd6916 : data_rom <= {16'd20169, 16'd25824};
                15'd6917 : data_rom <= {16'd20172, 16'd25822};
                15'd6918 : data_rom <= {16'd20174, 16'd25820};
                15'd6919 : data_rom <= {16'd20177, 16'd25819};
                15'd6920 : data_rom <= {16'd20179, 16'd25817};
                15'd6921 : data_rom <= {16'd20182, 16'd25815};
                15'd6922 : data_rom <= {16'd20184, 16'd25813};
                15'd6923 : data_rom <= {16'd20187, 16'd25811};
                15'd6924 : data_rom <= {16'd20189, 16'd25809};
                15'd6925 : data_rom <= {16'd20192, 16'd25807};
                15'd6926 : data_rom <= {16'd20194, 16'd25805};
                15'd6927 : data_rom <= {16'd20197, 16'd25803};
                15'd6928 : data_rom <= {16'd20199, 16'd25801};
                15'd6929 : data_rom <= {16'd20201, 16'd25799};
                15'd6930 : data_rom <= {16'd20204, 16'd25797};
                15'd6931 : data_rom <= {16'd20206, 16'd25795};
                15'd6932 : data_rom <= {16'd20209, 16'd25793};
                15'd6933 : data_rom <= {16'd20211, 16'd25791};
                15'd6934 : data_rom <= {16'd20214, 16'd25789};
                15'd6935 : data_rom <= {16'd20216, 16'd25788};
                15'd6936 : data_rom <= {16'd20219, 16'd25786};
                15'd6937 : data_rom <= {16'd20221, 16'd25784};
                15'd6938 : data_rom <= {16'd20224, 16'd25782};
                15'd6939 : data_rom <= {16'd20226, 16'd25780};
                15'd6940 : data_rom <= {16'd20229, 16'd25778};
                15'd6941 : data_rom <= {16'd20231, 16'd25776};
                15'd6942 : data_rom <= {16'd20234, 16'd25774};
                15'd6943 : data_rom <= {16'd20236, 16'd25772};
                15'd6944 : data_rom <= {16'd20239, 16'd25770};
                15'd6945 : data_rom <= {16'd20241, 16'd25768};
                15'd6946 : data_rom <= {16'd20243, 16'd25766};
                15'd6947 : data_rom <= {16'd20246, 16'd25764};
                15'd6948 : data_rom <= {16'd20248, 16'd25762};
                15'd6949 : data_rom <= {16'd20251, 16'd25760};
                15'd6950 : data_rom <= {16'd20253, 16'd25758};
                15'd6951 : data_rom <= {16'd20256, 16'd25756};
                15'd6952 : data_rom <= {16'd20258, 16'd25755};
                15'd6953 : data_rom <= {16'd20261, 16'd25753};
                15'd6954 : data_rom <= {16'd20263, 16'd25751};
                15'd6955 : data_rom <= {16'd20266, 16'd25749};
                15'd6956 : data_rom <= {16'd20268, 16'd25747};
                15'd6957 : data_rom <= {16'd20271, 16'd25745};
                15'd6958 : data_rom <= {16'd20273, 16'd25743};
                15'd6959 : data_rom <= {16'd20276, 16'd25741};
                15'd6960 : data_rom <= {16'd20278, 16'd25739};
                15'd6961 : data_rom <= {16'd20281, 16'd25737};
                15'd6962 : data_rom <= {16'd20283, 16'd25735};
                15'd6963 : data_rom <= {16'd20285, 16'd25733};
                15'd6964 : data_rom <= {16'd20288, 16'd25731};
                15'd6965 : data_rom <= {16'd20290, 16'd25729};
                15'd6966 : data_rom <= {16'd20293, 16'd25727};
                15'd6967 : data_rom <= {16'd20295, 16'd25725};
                15'd6968 : data_rom <= {16'd20298, 16'd25723};
                15'd6969 : data_rom <= {16'd20300, 16'd25721};
                15'd6970 : data_rom <= {16'd20303, 16'd25720};
                15'd6971 : data_rom <= {16'd20305, 16'd25718};
                15'd6972 : data_rom <= {16'd20308, 16'd25716};
                15'd6973 : data_rom <= {16'd20310, 16'd25714};
                15'd6974 : data_rom <= {16'd20313, 16'd25712};
                15'd6975 : data_rom <= {16'd20315, 16'd25710};
                15'd6976 : data_rom <= {16'd20318, 16'd25708};
                15'd6977 : data_rom <= {16'd20320, 16'd25706};
                15'd6978 : data_rom <= {16'd20322, 16'd25704};
                15'd6979 : data_rom <= {16'd20325, 16'd25702};
                15'd6980 : data_rom <= {16'd20327, 16'd25700};
                15'd6981 : data_rom <= {16'd20330, 16'd25698};
                15'd6982 : data_rom <= {16'd20332, 16'd25696};
                15'd6983 : data_rom <= {16'd20335, 16'd25694};
                15'd6984 : data_rom <= {16'd20337, 16'd25692};
                15'd6985 : data_rom <= {16'd20340, 16'd25690};
                15'd6986 : data_rom <= {16'd20342, 16'd25688};
                15'd6987 : data_rom <= {16'd20345, 16'd25686};
                15'd6988 : data_rom <= {16'd20347, 16'd25684};
                15'd6989 : data_rom <= {16'd20350, 16'd25683};
                15'd6990 : data_rom <= {16'd20352, 16'd25681};
                15'd6991 : data_rom <= {16'd20354, 16'd25679};
                15'd6992 : data_rom <= {16'd20357, 16'd25677};
                15'd6993 : data_rom <= {16'd20359, 16'd25675};
                15'd6994 : data_rom <= {16'd20362, 16'd25673};
                15'd6995 : data_rom <= {16'd20364, 16'd25671};
                15'd6996 : data_rom <= {16'd20367, 16'd25669};
                15'd6997 : data_rom <= {16'd20369, 16'd25667};
                15'd6998 : data_rom <= {16'd20372, 16'd25665};
                15'd6999 : data_rom <= {16'd20374, 16'd25663};
                15'd7000 : data_rom <= {16'd20377, 16'd25661};
                15'd7001 : data_rom <= {16'd20379, 16'd25659};
                15'd7002 : data_rom <= {16'd20382, 16'd25657};
                15'd7003 : data_rom <= {16'd20384, 16'd25655};
                15'd7004 : data_rom <= {16'd20386, 16'd25653};
                15'd7005 : data_rom <= {16'd20389, 16'd25651};
                15'd7006 : data_rom <= {16'd20391, 16'd25649};
                15'd7007 : data_rom <= {16'd20394, 16'd25647};
                15'd7008 : data_rom <= {16'd20396, 16'd25645};
                15'd7009 : data_rom <= {16'd20399, 16'd25643};
                15'd7010 : data_rom <= {16'd20401, 16'd25641};
                15'd7011 : data_rom <= {16'd20404, 16'd25640};
                15'd7012 : data_rom <= {16'd20406, 16'd25638};
                15'd7013 : data_rom <= {16'd20409, 16'd25636};
                15'd7014 : data_rom <= {16'd20411, 16'd25634};
                15'd7015 : data_rom <= {16'd20414, 16'd25632};
                15'd7016 : data_rom <= {16'd20416, 16'd25630};
                15'd7017 : data_rom <= {16'd20418, 16'd25628};
                15'd7018 : data_rom <= {16'd20421, 16'd25626};
                15'd7019 : data_rom <= {16'd20423, 16'd25624};
                15'd7020 : data_rom <= {16'd20426, 16'd25622};
                15'd7021 : data_rom <= {16'd20428, 16'd25620};
                15'd7022 : data_rom <= {16'd20431, 16'd25618};
                15'd7023 : data_rom <= {16'd20433, 16'd25616};
                15'd7024 : data_rom <= {16'd20436, 16'd25614};
                15'd7025 : data_rom <= {16'd20438, 16'd25612};
                15'd7026 : data_rom <= {16'd20441, 16'd25610};
                15'd7027 : data_rom <= {16'd20443, 16'd25608};
                15'd7028 : data_rom <= {16'd20445, 16'd25606};
                15'd7029 : data_rom <= {16'd20448, 16'd25604};
                15'd7030 : data_rom <= {16'd20450, 16'd25602};
                15'd7031 : data_rom <= {16'd20453, 16'd25600};
                15'd7032 : data_rom <= {16'd20455, 16'd25598};
                15'd7033 : data_rom <= {16'd20458, 16'd25596};
                15'd7034 : data_rom <= {16'd20460, 16'd25594};
                15'd7035 : data_rom <= {16'd20463, 16'd25593};
                15'd7036 : data_rom <= {16'd20465, 16'd25591};
                15'd7037 : data_rom <= {16'd20468, 16'd25589};
                15'd7038 : data_rom <= {16'd20470, 16'd25587};
                15'd7039 : data_rom <= {16'd20472, 16'd25585};
                15'd7040 : data_rom <= {16'd20475, 16'd25583};
                15'd7041 : data_rom <= {16'd20477, 16'd25581};
                15'd7042 : data_rom <= {16'd20480, 16'd25579};
                15'd7043 : data_rom <= {16'd20482, 16'd25577};
                15'd7044 : data_rom <= {16'd20485, 16'd25575};
                15'd7045 : data_rom <= {16'd20487, 16'd25573};
                15'd7046 : data_rom <= {16'd20490, 16'd25571};
                15'd7047 : data_rom <= {16'd20492, 16'd25569};
                15'd7048 : data_rom <= {16'd20494, 16'd25567};
                15'd7049 : data_rom <= {16'd20497, 16'd25565};
                15'd7050 : data_rom <= {16'd20499, 16'd25563};
                15'd7051 : data_rom <= {16'd20502, 16'd25561};
                15'd7052 : data_rom <= {16'd20504, 16'd25559};
                15'd7053 : data_rom <= {16'd20507, 16'd25557};
                15'd7054 : data_rom <= {16'd20509, 16'd25555};
                15'd7055 : data_rom <= {16'd20512, 16'd25553};
                15'd7056 : data_rom <= {16'd20514, 16'd25551};
                15'd7057 : data_rom <= {16'd20517, 16'd25549};
                15'd7058 : data_rom <= {16'd20519, 16'd25547};
                15'd7059 : data_rom <= {16'd20521, 16'd25545};
                15'd7060 : data_rom <= {16'd20524, 16'd25543};
                15'd7061 : data_rom <= {16'd20526, 16'd25541};
                15'd7062 : data_rom <= {16'd20529, 16'd25539};
                15'd7063 : data_rom <= {16'd20531, 16'd25537};
                15'd7064 : data_rom <= {16'd20534, 16'd25536};
                15'd7065 : data_rom <= {16'd20536, 16'd25534};
                15'd7066 : data_rom <= {16'd20539, 16'd25532};
                15'd7067 : data_rom <= {16'd20541, 16'd25530};
                15'd7068 : data_rom <= {16'd20543, 16'd25528};
                15'd7069 : data_rom <= {16'd20546, 16'd25526};
                15'd7070 : data_rom <= {16'd20548, 16'd25524};
                15'd7071 : data_rom <= {16'd20551, 16'd25522};
                15'd7072 : data_rom <= {16'd20553, 16'd25520};
                15'd7073 : data_rom <= {16'd20556, 16'd25518};
                15'd7074 : data_rom <= {16'd20558, 16'd25516};
                15'd7075 : data_rom <= {16'd20561, 16'd25514};
                15'd7076 : data_rom <= {16'd20563, 16'd25512};
                15'd7077 : data_rom <= {16'd20566, 16'd25510};
                15'd7078 : data_rom <= {16'd20568, 16'd25508};
                15'd7079 : data_rom <= {16'd20570, 16'd25506};
                15'd7080 : data_rom <= {16'd20573, 16'd25504};
                15'd7081 : data_rom <= {16'd20575, 16'd25502};
                15'd7082 : data_rom <= {16'd20578, 16'd25500};
                15'd7083 : data_rom <= {16'd20580, 16'd25498};
                15'd7084 : data_rom <= {16'd20583, 16'd25496};
                15'd7085 : data_rom <= {16'd20585, 16'd25494};
                15'd7086 : data_rom <= {16'd20588, 16'd25492};
                15'd7087 : data_rom <= {16'd20590, 16'd25490};
                15'd7088 : data_rom <= {16'd20592, 16'd25488};
                15'd7089 : data_rom <= {16'd20595, 16'd25486};
                15'd7090 : data_rom <= {16'd20597, 16'd25484};
                15'd7091 : data_rom <= {16'd20600, 16'd25482};
                15'd7092 : data_rom <= {16'd20602, 16'd25480};
                15'd7093 : data_rom <= {16'd20605, 16'd25478};
                15'd7094 : data_rom <= {16'd20607, 16'd25476};
                15'd7095 : data_rom <= {16'd20609, 16'd25474};
                15'd7096 : data_rom <= {16'd20612, 16'd25472};
                15'd7097 : data_rom <= {16'd20614, 16'd25470};
                15'd7098 : data_rom <= {16'd20617, 16'd25468};
                15'd7099 : data_rom <= {16'd20619, 16'd25466};
                15'd7100 : data_rom <= {16'd20622, 16'd25465};
                15'd7101 : data_rom <= {16'd20624, 16'd25463};
                15'd7102 : data_rom <= {16'd20627, 16'd25461};
                15'd7103 : data_rom <= {16'd20629, 16'd25459};
                15'd7104 : data_rom <= {16'd20631, 16'd25457};
                15'd7105 : data_rom <= {16'd20634, 16'd25455};
                15'd7106 : data_rom <= {16'd20636, 16'd25453};
                15'd7107 : data_rom <= {16'd20639, 16'd25451};
                15'd7108 : data_rom <= {16'd20641, 16'd25449};
                15'd7109 : data_rom <= {16'd20644, 16'd25447};
                15'd7110 : data_rom <= {16'd20646, 16'd25445};
                15'd7111 : data_rom <= {16'd20649, 16'd25443};
                15'd7112 : data_rom <= {16'd20651, 16'd25441};
                15'd7113 : data_rom <= {16'd20653, 16'd25439};
                15'd7114 : data_rom <= {16'd20656, 16'd25437};
                15'd7115 : data_rom <= {16'd20658, 16'd25435};
                15'd7116 : data_rom <= {16'd20661, 16'd25433};
                15'd7117 : data_rom <= {16'd20663, 16'd25431};
                15'd7118 : data_rom <= {16'd20666, 16'd25429};
                15'd7119 : data_rom <= {16'd20668, 16'd25427};
                15'd7120 : data_rom <= {16'd20670, 16'd25425};
                15'd7121 : data_rom <= {16'd20673, 16'd25423};
                15'd7122 : data_rom <= {16'd20675, 16'd25421};
                15'd7123 : data_rom <= {16'd20678, 16'd25419};
                15'd7124 : data_rom <= {16'd20680, 16'd25417};
                15'd7125 : data_rom <= {16'd20683, 16'd25415};
                15'd7126 : data_rom <= {16'd20685, 16'd25413};
                15'd7127 : data_rom <= {16'd20688, 16'd25411};
                15'd7128 : data_rom <= {16'd20690, 16'd25409};
                15'd7129 : data_rom <= {16'd20692, 16'd25407};
                15'd7130 : data_rom <= {16'd20695, 16'd25405};
                15'd7131 : data_rom <= {16'd20697, 16'd25403};
                15'd7132 : data_rom <= {16'd20700, 16'd25401};
                15'd7133 : data_rom <= {16'd20702, 16'd25399};
                15'd7134 : data_rom <= {16'd20705, 16'd25397};
                15'd7135 : data_rom <= {16'd20707, 16'd25395};
                15'd7136 : data_rom <= {16'd20709, 16'd25393};
                15'd7137 : data_rom <= {16'd20712, 16'd25391};
                15'd7138 : data_rom <= {16'd20714, 16'd25389};
                15'd7139 : data_rom <= {16'd20717, 16'd25387};
                15'd7140 : data_rom <= {16'd20719, 16'd25385};
                15'd7141 : data_rom <= {16'd20722, 16'd25383};
                15'd7142 : data_rom <= {16'd20724, 16'd25381};
                15'd7143 : data_rom <= {16'd20727, 16'd25379};
                15'd7144 : data_rom <= {16'd20729, 16'd25377};
                15'd7145 : data_rom <= {16'd20731, 16'd25375};
                15'd7146 : data_rom <= {16'd20734, 16'd25373};
                15'd7147 : data_rom <= {16'd20736, 16'd25371};
                15'd7148 : data_rom <= {16'd20739, 16'd25369};
                15'd7149 : data_rom <= {16'd20741, 16'd25367};
                15'd7150 : data_rom <= {16'd20744, 16'd25365};
                15'd7151 : data_rom <= {16'd20746, 16'd25363};
                15'd7152 : data_rom <= {16'd20748, 16'd25361};
                15'd7153 : data_rom <= {16'd20751, 16'd25359};
                15'd7154 : data_rom <= {16'd20753, 16'd25357};
                15'd7155 : data_rom <= {16'd20756, 16'd25355};
                15'd7156 : data_rom <= {16'd20758, 16'd25353};
                15'd7157 : data_rom <= {16'd20761, 16'd25351};
                15'd7158 : data_rom <= {16'd20763, 16'd25349};
                15'd7159 : data_rom <= {16'd20765, 16'd25347};
                15'd7160 : data_rom <= {16'd20768, 16'd25345};
                15'd7161 : data_rom <= {16'd20770, 16'd25343};
                15'd7162 : data_rom <= {16'd20773, 16'd25341};
                15'd7163 : data_rom <= {16'd20775, 16'd25339};
                15'd7164 : data_rom <= {16'd20778, 16'd25337};
                15'd7165 : data_rom <= {16'd20780, 16'd25335};
                15'd7166 : data_rom <= {16'd20782, 16'd25334};
                15'd7167 : data_rom <= {16'd20785, 16'd25332};
                15'd7168 : data_rom <= {16'd20787, 16'd25330};
                15'd7169 : data_rom <= {16'd20790, 16'd25328};
                15'd7170 : data_rom <= {16'd20792, 16'd25326};
                15'd7171 : data_rom <= {16'd20795, 16'd25324};
                15'd7172 : data_rom <= {16'd20797, 16'd25322};
                15'd7173 : data_rom <= {16'd20799, 16'd25320};
                15'd7174 : data_rom <= {16'd20802, 16'd25318};
                15'd7175 : data_rom <= {16'd20804, 16'd25316};
                15'd7176 : data_rom <= {16'd20807, 16'd25314};
                15'd7177 : data_rom <= {16'd20809, 16'd25312};
                15'd7178 : data_rom <= {16'd20812, 16'd25310};
                15'd7179 : data_rom <= {16'd20814, 16'd25308};
                15'd7180 : data_rom <= {16'd20816, 16'd25306};
                15'd7181 : data_rom <= {16'd20819, 16'd25304};
                15'd7182 : data_rom <= {16'd20821, 16'd25302};
                15'd7183 : data_rom <= {16'd20824, 16'd25300};
                15'd7184 : data_rom <= {16'd20826, 16'd25298};
                15'd7185 : data_rom <= {16'd20829, 16'd25296};
                15'd7186 : data_rom <= {16'd20831, 16'd25294};
                15'd7187 : data_rom <= {16'd20833, 16'd25292};
                15'd7188 : data_rom <= {16'd20836, 16'd25290};
                15'd7189 : data_rom <= {16'd20838, 16'd25288};
                15'd7190 : data_rom <= {16'd20841, 16'd25286};
                15'd7191 : data_rom <= {16'd20843, 16'd25284};
                15'd7192 : data_rom <= {16'd20846, 16'd25282};
                15'd7193 : data_rom <= {16'd20848, 16'd25280};
                15'd7194 : data_rom <= {16'd20850, 16'd25278};
                15'd7195 : data_rom <= {16'd20853, 16'd25276};
                15'd7196 : data_rom <= {16'd20855, 16'd25274};
                15'd7197 : data_rom <= {16'd20858, 16'd25272};
                15'd7198 : data_rom <= {16'd20860, 16'd25270};
                15'd7199 : data_rom <= {16'd20862, 16'd25268};
                15'd7200 : data_rom <= {16'd20865, 16'd25266};
                15'd7201 : data_rom <= {16'd20867, 16'd25264};
                15'd7202 : data_rom <= {16'd20870, 16'd25262};
                15'd7203 : data_rom <= {16'd20872, 16'd25260};
                15'd7204 : data_rom <= {16'd20875, 16'd25258};
                15'd7205 : data_rom <= {16'd20877, 16'd25256};
                15'd7206 : data_rom <= {16'd20879, 16'd25254};
                15'd7207 : data_rom <= {16'd20882, 16'd25252};
                15'd7208 : data_rom <= {16'd20884, 16'd25250};
                15'd7209 : data_rom <= {16'd20887, 16'd25248};
                15'd7210 : data_rom <= {16'd20889, 16'd25246};
                15'd7211 : data_rom <= {16'd20892, 16'd25244};
                15'd7212 : data_rom <= {16'd20894, 16'd25242};
                15'd7213 : data_rom <= {16'd20896, 16'd25240};
                15'd7214 : data_rom <= {16'd20899, 16'd25238};
                15'd7215 : data_rom <= {16'd20901, 16'd25236};
                15'd7216 : data_rom <= {16'd20904, 16'd25234};
                15'd7217 : data_rom <= {16'd20906, 16'd25232};
                15'd7218 : data_rom <= {16'd20908, 16'd25230};
                15'd7219 : data_rom <= {16'd20911, 16'd25228};
                15'd7220 : data_rom <= {16'd20913, 16'd25226};
                15'd7221 : data_rom <= {16'd20916, 16'd25224};
                15'd7222 : data_rom <= {16'd20918, 16'd25222};
                15'd7223 : data_rom <= {16'd20921, 16'd25220};
                15'd7224 : data_rom <= {16'd20923, 16'd25218};
                15'd7225 : data_rom <= {16'd20925, 16'd25216};
                15'd7226 : data_rom <= {16'd20928, 16'd25214};
                15'd7227 : data_rom <= {16'd20930, 16'd25212};
                15'd7228 : data_rom <= {16'd20933, 16'd25210};
                15'd7229 : data_rom <= {16'd20935, 16'd25208};
                15'd7230 : data_rom <= {16'd20937, 16'd25206};
                15'd7231 : data_rom <= {16'd20940, 16'd25203};
                15'd7232 : data_rom <= {16'd20942, 16'd25201};
                15'd7233 : data_rom <= {16'd20945, 16'd25199};
                15'd7234 : data_rom <= {16'd20947, 16'd25197};
                15'd7235 : data_rom <= {16'd20950, 16'd25195};
                15'd7236 : data_rom <= {16'd20952, 16'd25193};
                15'd7237 : data_rom <= {16'd20954, 16'd25191};
                15'd7238 : data_rom <= {16'd20957, 16'd25189};
                15'd7239 : data_rom <= {16'd20959, 16'd25187};
                15'd7240 : data_rom <= {16'd20962, 16'd25185};
                15'd7241 : data_rom <= {16'd20964, 16'd25183};
                15'd7242 : data_rom <= {16'd20966, 16'd25181};
                15'd7243 : data_rom <= {16'd20969, 16'd25179};
                15'd7244 : data_rom <= {16'd20971, 16'd25177};
                15'd7245 : data_rom <= {16'd20974, 16'd25175};
                15'd7246 : data_rom <= {16'd20976, 16'd25173};
                15'd7247 : data_rom <= {16'd20979, 16'd25171};
                15'd7248 : data_rom <= {16'd20981, 16'd25169};
                15'd7249 : data_rom <= {16'd20983, 16'd25167};
                15'd7250 : data_rom <= {16'd20986, 16'd25165};
                15'd7251 : data_rom <= {16'd20988, 16'd25163};
                15'd7252 : data_rom <= {16'd20991, 16'd25161};
                15'd7253 : data_rom <= {16'd20993, 16'd25159};
                15'd7254 : data_rom <= {16'd20995, 16'd25157};
                15'd7255 : data_rom <= {16'd20998, 16'd25155};
                15'd7256 : data_rom <= {16'd21000, 16'd25153};
                15'd7257 : data_rom <= {16'd21003, 16'd25151};
                15'd7258 : data_rom <= {16'd21005, 16'd25149};
                15'd7259 : data_rom <= {16'd21007, 16'd25147};
                15'd7260 : data_rom <= {16'd21010, 16'd25145};
                15'd7261 : data_rom <= {16'd21012, 16'd25143};
                15'd7262 : data_rom <= {16'd21015, 16'd25141};
                15'd7263 : data_rom <= {16'd21017, 16'd25139};
                15'd7264 : data_rom <= {16'd21020, 16'd25137};
                15'd7265 : data_rom <= {16'd21022, 16'd25135};
                15'd7266 : data_rom <= {16'd21024, 16'd25133};
                15'd7267 : data_rom <= {16'd21027, 16'd25131};
                15'd7268 : data_rom <= {16'd21029, 16'd25129};
                15'd7269 : data_rom <= {16'd21032, 16'd25127};
                15'd7270 : data_rom <= {16'd21034, 16'd25125};
                15'd7271 : data_rom <= {16'd21036, 16'd25123};
                15'd7272 : data_rom <= {16'd21039, 16'd25121};
                15'd7273 : data_rom <= {16'd21041, 16'd25119};
                15'd7274 : data_rom <= {16'd21044, 16'd25117};
                15'd7275 : data_rom <= {16'd21046, 16'd25115};
                15'd7276 : data_rom <= {16'd21048, 16'd25113};
                15'd7277 : data_rom <= {16'd21051, 16'd25111};
                15'd7278 : data_rom <= {16'd21053, 16'd25109};
                15'd7279 : data_rom <= {16'd21056, 16'd25107};
                15'd7280 : data_rom <= {16'd21058, 16'd25105};
                15'd7281 : data_rom <= {16'd21060, 16'd25103};
                15'd7282 : data_rom <= {16'd21063, 16'd25101};
                15'd7283 : data_rom <= {16'd21065, 16'd25099};
                15'd7284 : data_rom <= {16'd21068, 16'd25097};
                15'd7285 : data_rom <= {16'd21070, 16'd25095};
                15'd7286 : data_rom <= {16'd21073, 16'd25093};
                15'd7287 : data_rom <= {16'd21075, 16'd25091};
                15'd7288 : data_rom <= {16'd21077, 16'd25089};
                15'd7289 : data_rom <= {16'd21080, 16'd25087};
                15'd7290 : data_rom <= {16'd21082, 16'd25085};
                15'd7291 : data_rom <= {16'd21085, 16'd25083};
                15'd7292 : data_rom <= {16'd21087, 16'd25081};
                15'd7293 : data_rom <= {16'd21089, 16'd25079};
                15'd7294 : data_rom <= {16'd21092, 16'd25077};
                15'd7295 : data_rom <= {16'd21094, 16'd25075};
                15'd7296 : data_rom <= {16'd21097, 16'd25073};
                15'd7297 : data_rom <= {16'd21099, 16'd25070};
                15'd7298 : data_rom <= {16'd21101, 16'd25068};
                15'd7299 : data_rom <= {16'd21104, 16'd25066};
                15'd7300 : data_rom <= {16'd21106, 16'd25064};
                15'd7301 : data_rom <= {16'd21109, 16'd25062};
                15'd7302 : data_rom <= {16'd21111, 16'd25060};
                15'd7303 : data_rom <= {16'd21113, 16'd25058};
                15'd7304 : data_rom <= {16'd21116, 16'd25056};
                15'd7305 : data_rom <= {16'd21118, 16'd25054};
                15'd7306 : data_rom <= {16'd21121, 16'd25052};
                15'd7307 : data_rom <= {16'd21123, 16'd25050};
                15'd7308 : data_rom <= {16'd21125, 16'd25048};
                15'd7309 : data_rom <= {16'd21128, 16'd25046};
                15'd7310 : data_rom <= {16'd21130, 16'd25044};
                15'd7311 : data_rom <= {16'd21133, 16'd25042};
                15'd7312 : data_rom <= {16'd21135, 16'd25040};
                15'd7313 : data_rom <= {16'd21137, 16'd25038};
                15'd7314 : data_rom <= {16'd21140, 16'd25036};
                15'd7315 : data_rom <= {16'd21142, 16'd25034};
                15'd7316 : data_rom <= {16'd21145, 16'd25032};
                15'd7317 : data_rom <= {16'd21147, 16'd25030};
                15'd7318 : data_rom <= {16'd21149, 16'd25028};
                15'd7319 : data_rom <= {16'd21152, 16'd25026};
                15'd7320 : data_rom <= {16'd21154, 16'd25024};
                15'd7321 : data_rom <= {16'd21157, 16'd25022};
                15'd7322 : data_rom <= {16'd21159, 16'd25020};
                15'd7323 : data_rom <= {16'd21161, 16'd25018};
                15'd7324 : data_rom <= {16'd21164, 16'd25016};
                15'd7325 : data_rom <= {16'd21166, 16'd25014};
                15'd7326 : data_rom <= {16'd21169, 16'd25012};
                15'd7327 : data_rom <= {16'd21171, 16'd25010};
                15'd7328 : data_rom <= {16'd21173, 16'd25008};
                15'd7329 : data_rom <= {16'd21176, 16'd25006};
                15'd7330 : data_rom <= {16'd21178, 16'd25004};
                15'd7331 : data_rom <= {16'd21181, 16'd25002};
                15'd7332 : data_rom <= {16'd21183, 16'd25000};
                15'd7333 : data_rom <= {16'd21185, 16'd24998};
                15'd7334 : data_rom <= {16'd21188, 16'd24995};
                15'd7335 : data_rom <= {16'd21190, 16'd24993};
                15'd7336 : data_rom <= {16'd21193, 16'd24991};
                15'd7337 : data_rom <= {16'd21195, 16'd24989};
                15'd7338 : data_rom <= {16'd21197, 16'd24987};
                15'd7339 : data_rom <= {16'd21200, 16'd24985};
                15'd7340 : data_rom <= {16'd21202, 16'd24983};
                15'd7341 : data_rom <= {16'd21205, 16'd24981};
                15'd7342 : data_rom <= {16'd21207, 16'd24979};
                15'd7343 : data_rom <= {16'd21209, 16'd24977};
                15'd7344 : data_rom <= {16'd21212, 16'd24975};
                15'd7345 : data_rom <= {16'd21214, 16'd24973};
                15'd7346 : data_rom <= {16'd21217, 16'd24971};
                15'd7347 : data_rom <= {16'd21219, 16'd24969};
                15'd7348 : data_rom <= {16'd21221, 16'd24967};
                15'd7349 : data_rom <= {16'd21224, 16'd24965};
                15'd7350 : data_rom <= {16'd21226, 16'd24963};
                15'd7351 : data_rom <= {16'd21228, 16'd24961};
                15'd7352 : data_rom <= {16'd21231, 16'd24959};
                15'd7353 : data_rom <= {16'd21233, 16'd24957};
                15'd7354 : data_rom <= {16'd21236, 16'd24955};
                15'd7355 : data_rom <= {16'd21238, 16'd24953};
                15'd7356 : data_rom <= {16'd21240, 16'd24951};
                15'd7357 : data_rom <= {16'd21243, 16'd24949};
                15'd7358 : data_rom <= {16'd21245, 16'd24947};
                15'd7359 : data_rom <= {16'd21248, 16'd24945};
                15'd7360 : data_rom <= {16'd21250, 16'd24943};
                15'd7361 : data_rom <= {16'd21252, 16'd24941};
                15'd7362 : data_rom <= {16'd21255, 16'd24939};
                15'd7363 : data_rom <= {16'd21257, 16'd24936};
                15'd7364 : data_rom <= {16'd21260, 16'd24934};
                15'd7365 : data_rom <= {16'd21262, 16'd24932};
                15'd7366 : data_rom <= {16'd21264, 16'd24930};
                15'd7367 : data_rom <= {16'd21267, 16'd24928};
                15'd7368 : data_rom <= {16'd21269, 16'd24926};
                15'd7369 : data_rom <= {16'd21272, 16'd24924};
                15'd7370 : data_rom <= {16'd21274, 16'd24922};
                15'd7371 : data_rom <= {16'd21276, 16'd24920};
                15'd7372 : data_rom <= {16'd21279, 16'd24918};
                15'd7373 : data_rom <= {16'd21281, 16'd24916};
                15'd7374 : data_rom <= {16'd21283, 16'd24914};
                15'd7375 : data_rom <= {16'd21286, 16'd24912};
                15'd7376 : data_rom <= {16'd21288, 16'd24910};
                15'd7377 : data_rom <= {16'd21291, 16'd24908};
                15'd7378 : data_rom <= {16'd21293, 16'd24906};
                15'd7379 : data_rom <= {16'd21295, 16'd24904};
                15'd7380 : data_rom <= {16'd21298, 16'd24902};
                15'd7381 : data_rom <= {16'd21300, 16'd24900};
                15'd7382 : data_rom <= {16'd21303, 16'd24898};
                15'd7383 : data_rom <= {16'd21305, 16'd24896};
                15'd7384 : data_rom <= {16'd21307, 16'd24894};
                15'd7385 : data_rom <= {16'd21310, 16'd24892};
                15'd7386 : data_rom <= {16'd21312, 16'd24890};
                15'd7387 : data_rom <= {16'd21314, 16'd24888};
                15'd7388 : data_rom <= {16'd21317, 16'd24885};
                15'd7389 : data_rom <= {16'd21319, 16'd24883};
                15'd7390 : data_rom <= {16'd21322, 16'd24881};
                15'd7391 : data_rom <= {16'd21324, 16'd24879};
                15'd7392 : data_rom <= {16'd21326, 16'd24877};
                15'd7393 : data_rom <= {16'd21329, 16'd24875};
                15'd7394 : data_rom <= {16'd21331, 16'd24873};
                15'd7395 : data_rom <= {16'd21334, 16'd24871};
                15'd7396 : data_rom <= {16'd21336, 16'd24869};
                15'd7397 : data_rom <= {16'd21338, 16'd24867};
                15'd7398 : data_rom <= {16'd21341, 16'd24865};
                15'd7399 : data_rom <= {16'd21343, 16'd24863};
                15'd7400 : data_rom <= {16'd21346, 16'd24861};
                15'd7401 : data_rom <= {16'd21348, 16'd24859};
                15'd7402 : data_rom <= {16'd21350, 16'd24857};
                15'd7403 : data_rom <= {16'd21353, 16'd24855};
                15'd7404 : data_rom <= {16'd21355, 16'd24853};
                15'd7405 : data_rom <= {16'd21357, 16'd24851};
                15'd7406 : data_rom <= {16'd21360, 16'd24849};
                15'd7407 : data_rom <= {16'd21362, 16'd24847};
                15'd7408 : data_rom <= {16'd21365, 16'd24845};
                15'd7409 : data_rom <= {16'd21367, 16'd24842};
                15'd7410 : data_rom <= {16'd21369, 16'd24840};
                15'd7411 : data_rom <= {16'd21372, 16'd24838};
                15'd7412 : data_rom <= {16'd21374, 16'd24836};
                15'd7413 : data_rom <= {16'd21376, 16'd24834};
                15'd7414 : data_rom <= {16'd21379, 16'd24832};
                15'd7415 : data_rom <= {16'd21381, 16'd24830};
                15'd7416 : data_rom <= {16'd21384, 16'd24828};
                15'd7417 : data_rom <= {16'd21386, 16'd24826};
                15'd7418 : data_rom <= {16'd21388, 16'd24824};
                15'd7419 : data_rom <= {16'd21391, 16'd24822};
                15'd7420 : data_rom <= {16'd21393, 16'd24820};
                15'd7421 : data_rom <= {16'd21396, 16'd24818};
                15'd7422 : data_rom <= {16'd21398, 16'd24816};
                15'd7423 : data_rom <= {16'd21400, 16'd24814};
                15'd7424 : data_rom <= {16'd21403, 16'd24812};
                15'd7425 : data_rom <= {16'd21405, 16'd24810};
                15'd7426 : data_rom <= {16'd21407, 16'd24808};
                15'd7427 : data_rom <= {16'd21410, 16'd24806};
                15'd7428 : data_rom <= {16'd21412, 16'd24804};
                15'd7429 : data_rom <= {16'd21415, 16'd24801};
                15'd7430 : data_rom <= {16'd21417, 16'd24799};
                15'd7431 : data_rom <= {16'd21419, 16'd24797};
                15'd7432 : data_rom <= {16'd21422, 16'd24795};
                15'd7433 : data_rom <= {16'd21424, 16'd24793};
                15'd7434 : data_rom <= {16'd21426, 16'd24791};
                15'd7435 : data_rom <= {16'd21429, 16'd24789};
                15'd7436 : data_rom <= {16'd21431, 16'd24787};
                15'd7437 : data_rom <= {16'd21434, 16'd24785};
                15'd7438 : data_rom <= {16'd21436, 16'd24783};
                15'd7439 : data_rom <= {16'd21438, 16'd24781};
                15'd7440 : data_rom <= {16'd21441, 16'd24779};
                15'd7441 : data_rom <= {16'd21443, 16'd24777};
                15'd7442 : data_rom <= {16'd21445, 16'd24775};
                15'd7443 : data_rom <= {16'd21448, 16'd24773};
                15'd7444 : data_rom <= {16'd21450, 16'd24771};
                15'd7445 : data_rom <= {16'd21453, 16'd24769};
                15'd7446 : data_rom <= {16'd21455, 16'd24767};
                15'd7447 : data_rom <= {16'd21457, 16'd24764};
                15'd7448 : data_rom <= {16'd21460, 16'd24762};
                15'd7449 : data_rom <= {16'd21462, 16'd24760};
                15'd7450 : data_rom <= {16'd21464, 16'd24758};
                15'd7451 : data_rom <= {16'd21467, 16'd24756};
                15'd7452 : data_rom <= {16'd21469, 16'd24754};
                15'd7453 : data_rom <= {16'd21472, 16'd24752};
                15'd7454 : data_rom <= {16'd21474, 16'd24750};
                15'd7455 : data_rom <= {16'd21476, 16'd24748};
                15'd7456 : data_rom <= {16'd21479, 16'd24746};
                15'd7457 : data_rom <= {16'd21481, 16'd24744};
                15'd7458 : data_rom <= {16'd21483, 16'd24742};
                15'd7459 : data_rom <= {16'd21486, 16'd24740};
                15'd7460 : data_rom <= {16'd21488, 16'd24738};
                15'd7461 : data_rom <= {16'd21491, 16'd24736};
                15'd7462 : data_rom <= {16'd21493, 16'd24734};
                15'd7463 : data_rom <= {16'd21495, 16'd24732};
                15'd7464 : data_rom <= {16'd21498, 16'd24729};
                15'd7465 : data_rom <= {16'd21500, 16'd24727};
                15'd7466 : data_rom <= {16'd21502, 16'd24725};
                15'd7467 : data_rom <= {16'd21505, 16'd24723};
                15'd7468 : data_rom <= {16'd21507, 16'd24721};
                15'd7469 : data_rom <= {16'd21509, 16'd24719};
                15'd7470 : data_rom <= {16'd21512, 16'd24717};
                15'd7471 : data_rom <= {16'd21514, 16'd24715};
                15'd7472 : data_rom <= {16'd21517, 16'd24713};
                15'd7473 : data_rom <= {16'd21519, 16'd24711};
                15'd7474 : data_rom <= {16'd21521, 16'd24709};
                15'd7475 : data_rom <= {16'd21524, 16'd24707};
                15'd7476 : data_rom <= {16'd21526, 16'd24705};
                15'd7477 : data_rom <= {16'd21528, 16'd24703};
                15'd7478 : data_rom <= {16'd21531, 16'd24701};
                15'd7479 : data_rom <= {16'd21533, 16'd24699};
                15'd7480 : data_rom <= {16'd21536, 16'd24696};
                15'd7481 : data_rom <= {16'd21538, 16'd24694};
                15'd7482 : data_rom <= {16'd21540, 16'd24692};
                15'd7483 : data_rom <= {16'd21543, 16'd24690};
                15'd7484 : data_rom <= {16'd21545, 16'd24688};
                15'd7485 : data_rom <= {16'd21547, 16'd24686};
                15'd7486 : data_rom <= {16'd21550, 16'd24684};
                15'd7487 : data_rom <= {16'd21552, 16'd24682};
                15'd7488 : data_rom <= {16'd21554, 16'd24680};
                15'd7489 : data_rom <= {16'd21557, 16'd24678};
                15'd7490 : data_rom <= {16'd21559, 16'd24676};
                15'd7491 : data_rom <= {16'd21562, 16'd24674};
                15'd7492 : data_rom <= {16'd21564, 16'd24672};
                15'd7493 : data_rom <= {16'd21566, 16'd24670};
                15'd7494 : data_rom <= {16'd21569, 16'd24668};
                15'd7495 : data_rom <= {16'd21571, 16'd24665};
                15'd7496 : data_rom <= {16'd21573, 16'd24663};
                15'd7497 : data_rom <= {16'd21576, 16'd24661};
                15'd7498 : data_rom <= {16'd21578, 16'd24659};
                15'd7499 : data_rom <= {16'd21581, 16'd24657};
                15'd7500 : data_rom <= {16'd21583, 16'd24655};
                15'd7501 : data_rom <= {16'd21585, 16'd24653};
                15'd7502 : data_rom <= {16'd21588, 16'd24651};
                15'd7503 : data_rom <= {16'd21590, 16'd24649};
                15'd7504 : data_rom <= {16'd21592, 16'd24647};
                15'd7505 : data_rom <= {16'd21595, 16'd24645};
                15'd7506 : data_rom <= {16'd21597, 16'd24643};
                15'd7507 : data_rom <= {16'd21599, 16'd24641};
                15'd7508 : data_rom <= {16'd21602, 16'd24639};
                15'd7509 : data_rom <= {16'd21604, 16'd24636};
                15'd7510 : data_rom <= {16'd21607, 16'd24634};
                15'd7511 : data_rom <= {16'd21609, 16'd24632};
                15'd7512 : data_rom <= {16'd21611, 16'd24630};
                15'd7513 : data_rom <= {16'd21614, 16'd24628};
                15'd7514 : data_rom <= {16'd21616, 16'd24626};
                15'd7515 : data_rom <= {16'd21618, 16'd24624};
                15'd7516 : data_rom <= {16'd21621, 16'd24622};
                15'd7517 : data_rom <= {16'd21623, 16'd24620};
                15'd7518 : data_rom <= {16'd21625, 16'd24618};
                15'd7519 : data_rom <= {16'd21628, 16'd24616};
                15'd7520 : data_rom <= {16'd21630, 16'd24614};
                15'd7521 : data_rom <= {16'd21632, 16'd24612};
                15'd7522 : data_rom <= {16'd21635, 16'd24610};
                15'd7523 : data_rom <= {16'd21637, 16'd24607};
                15'd7524 : data_rom <= {16'd21640, 16'd24605};
                15'd7525 : data_rom <= {16'd21642, 16'd24603};
                15'd7526 : data_rom <= {16'd21644, 16'd24601};
                15'd7527 : data_rom <= {16'd21647, 16'd24599};
                15'd7528 : data_rom <= {16'd21649, 16'd24597};
                15'd7529 : data_rom <= {16'd21651, 16'd24595};
                15'd7530 : data_rom <= {16'd21654, 16'd24593};
                15'd7531 : data_rom <= {16'd21656, 16'd24591};
                15'd7532 : data_rom <= {16'd21658, 16'd24589};
                15'd7533 : data_rom <= {16'd21661, 16'd24587};
                15'd7534 : data_rom <= {16'd21663, 16'd24585};
                15'd7535 : data_rom <= {16'd21665, 16'd24583};
                15'd7536 : data_rom <= {16'd21668, 16'd24580};
                15'd7537 : data_rom <= {16'd21670, 16'd24578};
                15'd7538 : data_rom <= {16'd21673, 16'd24576};
                15'd7539 : data_rom <= {16'd21675, 16'd24574};
                15'd7540 : data_rom <= {16'd21677, 16'd24572};
                15'd7541 : data_rom <= {16'd21680, 16'd24570};
                15'd7542 : data_rom <= {16'd21682, 16'd24568};
                15'd7543 : data_rom <= {16'd21684, 16'd24566};
                15'd7544 : data_rom <= {16'd21687, 16'd24564};
                15'd7545 : data_rom <= {16'd21689, 16'd24562};
                15'd7546 : data_rom <= {16'd21691, 16'd24560};
                15'd7547 : data_rom <= {16'd21694, 16'd24558};
                15'd7548 : data_rom <= {16'd21696, 16'd24556};
                15'd7549 : data_rom <= {16'd21698, 16'd24553};
                15'd7550 : data_rom <= {16'd21701, 16'd24551};
                15'd7551 : data_rom <= {16'd21703, 16'd24549};
                15'd7552 : data_rom <= {16'd21706, 16'd24547};
                15'd7553 : data_rom <= {16'd21708, 16'd24545};
                15'd7554 : data_rom <= {16'd21710, 16'd24543};
                15'd7555 : data_rom <= {16'd21713, 16'd24541};
                15'd7556 : data_rom <= {16'd21715, 16'd24539};
                15'd7557 : data_rom <= {16'd21717, 16'd24537};
                15'd7558 : data_rom <= {16'd21720, 16'd24535};
                15'd7559 : data_rom <= {16'd21722, 16'd24533};
                15'd7560 : data_rom <= {16'd21724, 16'd24531};
                15'd7561 : data_rom <= {16'd21727, 16'd24528};
                15'd7562 : data_rom <= {16'd21729, 16'd24526};
                15'd7563 : data_rom <= {16'd21731, 16'd24524};
                15'd7564 : data_rom <= {16'd21734, 16'd24522};
                15'd7565 : data_rom <= {16'd21736, 16'd24520};
                15'd7566 : data_rom <= {16'd21738, 16'd24518};
                15'd7567 : data_rom <= {16'd21741, 16'd24516};
                15'd7568 : data_rom <= {16'd21743, 16'd24514};
                15'd7569 : data_rom <= {16'd21746, 16'd24512};
                15'd7570 : data_rom <= {16'd21748, 16'd24510};
                15'd7571 : data_rom <= {16'd21750, 16'd24508};
                15'd7572 : data_rom <= {16'd21753, 16'd24506};
                15'd7573 : data_rom <= {16'd21755, 16'd24503};
                15'd7574 : data_rom <= {16'd21757, 16'd24501};
                15'd7575 : data_rom <= {16'd21760, 16'd24499};
                15'd7576 : data_rom <= {16'd21762, 16'd24497};
                15'd7577 : data_rom <= {16'd21764, 16'd24495};
                15'd7578 : data_rom <= {16'd21767, 16'd24493};
                15'd7579 : data_rom <= {16'd21769, 16'd24491};
                15'd7580 : data_rom <= {16'd21771, 16'd24489};
                15'd7581 : data_rom <= {16'd21774, 16'd24487};
                15'd7582 : data_rom <= {16'd21776, 16'd24485};
                15'd7583 : data_rom <= {16'd21778, 16'd24483};
                15'd7584 : data_rom <= {16'd21781, 16'd24481};
                15'd7585 : data_rom <= {16'd21783, 16'd24478};
                15'd7586 : data_rom <= {16'd21785, 16'd24476};
                15'd7587 : data_rom <= {16'd21788, 16'd24474};
                15'd7588 : data_rom <= {16'd21790, 16'd24472};
                15'd7589 : data_rom <= {16'd21792, 16'd24470};
                15'd7590 : data_rom <= {16'd21795, 16'd24468};
                15'd7591 : data_rom <= {16'd21797, 16'd24466};
                15'd7592 : data_rom <= {16'd21800, 16'd24464};
                15'd7593 : data_rom <= {16'd21802, 16'd24462};
                15'd7594 : data_rom <= {16'd21804, 16'd24460};
                15'd7595 : data_rom <= {16'd21807, 16'd24458};
                15'd7596 : data_rom <= {16'd21809, 16'd24455};
                15'd7597 : data_rom <= {16'd21811, 16'd24453};
                15'd7598 : data_rom <= {16'd21814, 16'd24451};
                15'd7599 : data_rom <= {16'd21816, 16'd24449};
                15'd7600 : data_rom <= {16'd21818, 16'd24447};
                15'd7601 : data_rom <= {16'd21821, 16'd24445};
                15'd7602 : data_rom <= {16'd21823, 16'd24443};
                15'd7603 : data_rom <= {16'd21825, 16'd24441};
                15'd7604 : data_rom <= {16'd21828, 16'd24439};
                15'd7605 : data_rom <= {16'd21830, 16'd24437};
                15'd7606 : data_rom <= {16'd21832, 16'd24435};
                15'd7607 : data_rom <= {16'd21835, 16'd24432};
                15'd7608 : data_rom <= {16'd21837, 16'd24430};
                15'd7609 : data_rom <= {16'd21839, 16'd24428};
                15'd7610 : data_rom <= {16'd21842, 16'd24426};
                15'd7611 : data_rom <= {16'd21844, 16'd24424};
                15'd7612 : data_rom <= {16'd21846, 16'd24422};
                15'd7613 : data_rom <= {16'd21849, 16'd24420};
                15'd7614 : data_rom <= {16'd21851, 16'd24418};
                15'd7615 : data_rom <= {16'd21853, 16'd24416};
                15'd7616 : data_rom <= {16'd21856, 16'd24414};
                15'd7617 : data_rom <= {16'd21858, 16'd24411};
                15'd7618 : data_rom <= {16'd21860, 16'd24409};
                15'd7619 : data_rom <= {16'd21863, 16'd24407};
                15'd7620 : data_rom <= {16'd21865, 16'd24405};
                15'd7621 : data_rom <= {16'd21867, 16'd24403};
                15'd7622 : data_rom <= {16'd21870, 16'd24401};
                15'd7623 : data_rom <= {16'd21872, 16'd24399};
                15'd7624 : data_rom <= {16'd21874, 16'd24397};
                15'd7625 : data_rom <= {16'd21877, 16'd24395};
                15'd7626 : data_rom <= {16'd21879, 16'd24393};
                15'd7627 : data_rom <= {16'd21881, 16'd24391};
                15'd7628 : data_rom <= {16'd21884, 16'd24388};
                15'd7629 : data_rom <= {16'd21886, 16'd24386};
                15'd7630 : data_rom <= {16'd21888, 16'd24384};
                15'd7631 : data_rom <= {16'd21891, 16'd24382};
                15'd7632 : data_rom <= {16'd21893, 16'd24380};
                15'd7633 : data_rom <= {16'd21895, 16'd24378};
                15'd7634 : data_rom <= {16'd21898, 16'd24376};
                15'd7635 : data_rom <= {16'd21900, 16'd24374};
                15'd7636 : data_rom <= {16'd21903, 16'd24372};
                15'd7637 : data_rom <= {16'd21905, 16'd24370};
                15'd7638 : data_rom <= {16'd21907, 16'd24367};
                15'd7639 : data_rom <= {16'd21910, 16'd24365};
                15'd7640 : data_rom <= {16'd21912, 16'd24363};
                15'd7641 : data_rom <= {16'd21914, 16'd24361};
                15'd7642 : data_rom <= {16'd21917, 16'd24359};
                15'd7643 : data_rom <= {16'd21919, 16'd24357};
                15'd7644 : data_rom <= {16'd21921, 16'd24355};
                15'd7645 : data_rom <= {16'd21924, 16'd24353};
                15'd7646 : data_rom <= {16'd21926, 16'd24351};
                15'd7647 : data_rom <= {16'd21928, 16'd24349};
                15'd7648 : data_rom <= {16'd21931, 16'd24346};
                15'd7649 : data_rom <= {16'd21933, 16'd24344};
                15'd7650 : data_rom <= {16'd21935, 16'd24342};
                15'd7651 : data_rom <= {16'd21938, 16'd24340};
                15'd7652 : data_rom <= {16'd21940, 16'd24338};
                15'd7653 : data_rom <= {16'd21942, 16'd24336};
                15'd7654 : data_rom <= {16'd21945, 16'd24334};
                15'd7655 : data_rom <= {16'd21947, 16'd24332};
                15'd7656 : data_rom <= {16'd21949, 16'd24330};
                15'd7657 : data_rom <= {16'd21952, 16'd24327};
                15'd7658 : data_rom <= {16'd21954, 16'd24325};
                15'd7659 : data_rom <= {16'd21956, 16'd24323};
                15'd7660 : data_rom <= {16'd21959, 16'd24321};
                15'd7661 : data_rom <= {16'd21961, 16'd24319};
                15'd7662 : data_rom <= {16'd21963, 16'd24317};
                15'd7663 : data_rom <= {16'd21966, 16'd24315};
                15'd7664 : data_rom <= {16'd21968, 16'd24313};
                15'd7665 : data_rom <= {16'd21970, 16'd24311};
                15'd7666 : data_rom <= {16'd21973, 16'd24309};
                15'd7667 : data_rom <= {16'd21975, 16'd24306};
                15'd7668 : data_rom <= {16'd21977, 16'd24304};
                15'd7669 : data_rom <= {16'd21980, 16'd24302};
                15'd7670 : data_rom <= {16'd21982, 16'd24300};
                15'd7671 : data_rom <= {16'd21984, 16'd24298};
                15'd7672 : data_rom <= {16'd21986, 16'd24296};
                15'd7673 : data_rom <= {16'd21989, 16'd24294};
                15'd7674 : data_rom <= {16'd21991, 16'd24292};
                15'd7675 : data_rom <= {16'd21993, 16'd24290};
                15'd7676 : data_rom <= {16'd21996, 16'd24287};
                15'd7677 : data_rom <= {16'd21998, 16'd24285};
                15'd7678 : data_rom <= {16'd22000, 16'd24283};
                15'd7679 : data_rom <= {16'd22003, 16'd24281};
                15'd7680 : data_rom <= {16'd22005, 16'd24279};
                15'd7681 : data_rom <= {16'd22007, 16'd24277};
                15'd7682 : data_rom <= {16'd22010, 16'd24275};
                15'd7683 : data_rom <= {16'd22012, 16'd24273};
                15'd7684 : data_rom <= {16'd22014, 16'd24271};
                15'd7685 : data_rom <= {16'd22017, 16'd24268};
                15'd7686 : data_rom <= {16'd22019, 16'd24266};
                15'd7687 : data_rom <= {16'd22021, 16'd24264};
                15'd7688 : data_rom <= {16'd22024, 16'd24262};
                15'd7689 : data_rom <= {16'd22026, 16'd24260};
                15'd7690 : data_rom <= {16'd22028, 16'd24258};
                15'd7691 : data_rom <= {16'd22031, 16'd24256};
                15'd7692 : data_rom <= {16'd22033, 16'd24254};
                15'd7693 : data_rom <= {16'd22035, 16'd24252};
                15'd7694 : data_rom <= {16'd22038, 16'd24249};
                15'd7695 : data_rom <= {16'd22040, 16'd24247};
                15'd7696 : data_rom <= {16'd22042, 16'd24245};
                15'd7697 : data_rom <= {16'd22045, 16'd24243};
                15'd7698 : data_rom <= {16'd22047, 16'd24241};
                15'd7699 : data_rom <= {16'd22049, 16'd24239};
                15'd7700 : data_rom <= {16'd22052, 16'd24237};
                15'd7701 : data_rom <= {16'd22054, 16'd24235};
                15'd7702 : data_rom <= {16'd22056, 16'd24233};
                15'd7703 : data_rom <= {16'd22059, 16'd24230};
                15'd7704 : data_rom <= {16'd22061, 16'd24228};
                15'd7705 : data_rom <= {16'd22063, 16'd24226};
                15'd7706 : data_rom <= {16'd22066, 16'd24224};
                15'd7707 : data_rom <= {16'd22068, 16'd24222};
                15'd7708 : data_rom <= {16'd22070, 16'd24220};
                15'd7709 : data_rom <= {16'd22073, 16'd24218};
                15'd7710 : data_rom <= {16'd22075, 16'd24216};
                15'd7711 : data_rom <= {16'd22077, 16'd24213};
                15'd7712 : data_rom <= {16'd22080, 16'd24211};
                15'd7713 : data_rom <= {16'd22082, 16'd24209};
                15'd7714 : data_rom <= {16'd22084, 16'd24207};
                15'd7715 : data_rom <= {16'd22086, 16'd24205};
                15'd7716 : data_rom <= {16'd22089, 16'd24203};
                15'd7717 : data_rom <= {16'd22091, 16'd24201};
                15'd7718 : data_rom <= {16'd22093, 16'd24199};
                15'd7719 : data_rom <= {16'd22096, 16'd24197};
                15'd7720 : data_rom <= {16'd22098, 16'd24194};
                15'd7721 : data_rom <= {16'd22100, 16'd24192};
                15'd7722 : data_rom <= {16'd22103, 16'd24190};
                15'd7723 : data_rom <= {16'd22105, 16'd24188};
                15'd7724 : data_rom <= {16'd22107, 16'd24186};
                15'd7725 : data_rom <= {16'd22110, 16'd24184};
                15'd7726 : data_rom <= {16'd22112, 16'd24182};
                15'd7727 : data_rom <= {16'd22114, 16'd24180};
                15'd7728 : data_rom <= {16'd22117, 16'd24177};
                15'd7729 : data_rom <= {16'd22119, 16'd24175};
                15'd7730 : data_rom <= {16'd22121, 16'd24173};
                15'd7731 : data_rom <= {16'd22124, 16'd24171};
                15'd7732 : data_rom <= {16'd22126, 16'd24169};
                15'd7733 : data_rom <= {16'd22128, 16'd24167};
                15'd7734 : data_rom <= {16'd22131, 16'd24165};
                15'd7735 : data_rom <= {16'd22133, 16'd24163};
                15'd7736 : data_rom <= {16'd22135, 16'd24161};
                15'd7737 : data_rom <= {16'd22137, 16'd24158};
                15'd7738 : data_rom <= {16'd22140, 16'd24156};
                15'd7739 : data_rom <= {16'd22142, 16'd24154};
                15'd7740 : data_rom <= {16'd22144, 16'd24152};
                15'd7741 : data_rom <= {16'd22147, 16'd24150};
                15'd7742 : data_rom <= {16'd22149, 16'd24148};
                15'd7743 : data_rom <= {16'd22151, 16'd24146};
                15'd7744 : data_rom <= {16'd22154, 16'd24144};
                15'd7745 : data_rom <= {16'd22156, 16'd24141};
                15'd7746 : data_rom <= {16'd22158, 16'd24139};
                15'd7747 : data_rom <= {16'd22161, 16'd24137};
                15'd7748 : data_rom <= {16'd22163, 16'd24135};
                15'd7749 : data_rom <= {16'd22165, 16'd24133};
                15'd7750 : data_rom <= {16'd22168, 16'd24131};
                15'd7751 : data_rom <= {16'd22170, 16'd24129};
                15'd7752 : data_rom <= {16'd22172, 16'd24127};
                15'd7753 : data_rom <= {16'd22175, 16'd24124};
                15'd7754 : data_rom <= {16'd22177, 16'd24122};
                15'd7755 : data_rom <= {16'd22179, 16'd24120};
                15'd7756 : data_rom <= {16'd22181, 16'd24118};
                15'd7757 : data_rom <= {16'd22184, 16'd24116};
                15'd7758 : data_rom <= {16'd22186, 16'd24114};
                15'd7759 : data_rom <= {16'd22188, 16'd24112};
                15'd7760 : data_rom <= {16'd22191, 16'd24110};
                15'd7761 : data_rom <= {16'd22193, 16'd24107};
                15'd7762 : data_rom <= {16'd22195, 16'd24105};
                15'd7763 : data_rom <= {16'd22198, 16'd24103};
                15'd7764 : data_rom <= {16'd22200, 16'd24101};
                15'd7765 : data_rom <= {16'd22202, 16'd24099};
                15'd7766 : data_rom <= {16'd22205, 16'd24097};
                15'd7767 : data_rom <= {16'd22207, 16'd24095};
                15'd7768 : data_rom <= {16'd22209, 16'd24092};
                15'd7769 : data_rom <= {16'd22211, 16'd24090};
                15'd7770 : data_rom <= {16'd22214, 16'd24088};
                15'd7771 : data_rom <= {16'd22216, 16'd24086};
                15'd7772 : data_rom <= {16'd22218, 16'd24084};
                15'd7773 : data_rom <= {16'd22221, 16'd24082};
                15'd7774 : data_rom <= {16'd22223, 16'd24080};
                15'd7775 : data_rom <= {16'd22225, 16'd24078};
                15'd7776 : data_rom <= {16'd22228, 16'd24075};
                15'd7777 : data_rom <= {16'd22230, 16'd24073};
                15'd7778 : data_rom <= {16'd22232, 16'd24071};
                15'd7779 : data_rom <= {16'd22235, 16'd24069};
                15'd7780 : data_rom <= {16'd22237, 16'd24067};
                15'd7781 : data_rom <= {16'd22239, 16'd24065};
                15'd7782 : data_rom <= {16'd22242, 16'd24063};
                15'd7783 : data_rom <= {16'd22244, 16'd24061};
                15'd7784 : data_rom <= {16'd22246, 16'd24058};
                15'd7785 : data_rom <= {16'd22248, 16'd24056};
                15'd7786 : data_rom <= {16'd22251, 16'd24054};
                15'd7787 : data_rom <= {16'd22253, 16'd24052};
                15'd7788 : data_rom <= {16'd22255, 16'd24050};
                15'd7789 : data_rom <= {16'd22258, 16'd24048};
                15'd7790 : data_rom <= {16'd22260, 16'd24046};
                15'd7791 : data_rom <= {16'd22262, 16'd24043};
                15'd7792 : data_rom <= {16'd22265, 16'd24041};
                15'd7793 : data_rom <= {16'd22267, 16'd24039};
                15'd7794 : data_rom <= {16'd22269, 16'd24037};
                15'd7795 : data_rom <= {16'd22271, 16'd24035};
                15'd7796 : data_rom <= {16'd22274, 16'd24033};
                15'd7797 : data_rom <= {16'd22276, 16'd24031};
                15'd7798 : data_rom <= {16'd22278, 16'd24029};
                15'd7799 : data_rom <= {16'd22281, 16'd24026};
                15'd7800 : data_rom <= {16'd22283, 16'd24024};
                15'd7801 : data_rom <= {16'd22285, 16'd24022};
                15'd7802 : data_rom <= {16'd22288, 16'd24020};
                15'd7803 : data_rom <= {16'd22290, 16'd24018};
                15'd7804 : data_rom <= {16'd22292, 16'd24016};
                15'd7805 : data_rom <= {16'd22295, 16'd24014};
                15'd7806 : data_rom <= {16'd22297, 16'd24011};
                15'd7807 : data_rom <= {16'd22299, 16'd24009};
                15'd7808 : data_rom <= {16'd22301, 16'd24007};
                15'd7809 : data_rom <= {16'd22304, 16'd24005};
                15'd7810 : data_rom <= {16'd22306, 16'd24003};
                15'd7811 : data_rom <= {16'd22308, 16'd24001};
                15'd7812 : data_rom <= {16'd22311, 16'd23999};
                15'd7813 : data_rom <= {16'd22313, 16'd23996};
                15'd7814 : data_rom <= {16'd22315, 16'd23994};
                15'd7815 : data_rom <= {16'd22318, 16'd23992};
                15'd7816 : data_rom <= {16'd22320, 16'd23990};
                15'd7817 : data_rom <= {16'd22322, 16'd23988};
                15'd7818 : data_rom <= {16'd22324, 16'd23986};
                15'd7819 : data_rom <= {16'd22327, 16'd23984};
                15'd7820 : data_rom <= {16'd22329, 16'd23981};
                15'd7821 : data_rom <= {16'd22331, 16'd23979};
                15'd7822 : data_rom <= {16'd22334, 16'd23977};
                15'd7823 : data_rom <= {16'd22336, 16'd23975};
                15'd7824 : data_rom <= {16'd22338, 16'd23973};
                15'd7825 : data_rom <= {16'd22341, 16'd23971};
                15'd7826 : data_rom <= {16'd22343, 16'd23969};
                15'd7827 : data_rom <= {16'd22345, 16'd23966};
                15'd7828 : data_rom <= {16'd22347, 16'd23964};
                15'd7829 : data_rom <= {16'd22350, 16'd23962};
                15'd7830 : data_rom <= {16'd22352, 16'd23960};
                15'd7831 : data_rom <= {16'd22354, 16'd23958};
                15'd7832 : data_rom <= {16'd22357, 16'd23956};
                15'd7833 : data_rom <= {16'd22359, 16'd23954};
                15'd7834 : data_rom <= {16'd22361, 16'd23951};
                15'd7835 : data_rom <= {16'd22363, 16'd23949};
                15'd7836 : data_rom <= {16'd22366, 16'd23947};
                15'd7837 : data_rom <= {16'd22368, 16'd23945};
                15'd7838 : data_rom <= {16'd22370, 16'd23943};
                15'd7839 : data_rom <= {16'd22373, 16'd23941};
                15'd7840 : data_rom <= {16'd22375, 16'd23939};
                15'd7841 : data_rom <= {16'd22377, 16'd23936};
                15'd7842 : data_rom <= {16'd22380, 16'd23934};
                15'd7843 : data_rom <= {16'd22382, 16'd23932};
                15'd7844 : data_rom <= {16'd22384, 16'd23930};
                15'd7845 : data_rom <= {16'd22386, 16'd23928};
                15'd7846 : data_rom <= {16'd22389, 16'd23926};
                15'd7847 : data_rom <= {16'd22391, 16'd23924};
                15'd7848 : data_rom <= {16'd22393, 16'd23921};
                15'd7849 : data_rom <= {16'd22396, 16'd23919};
                15'd7850 : data_rom <= {16'd22398, 16'd23917};
                15'd7851 : data_rom <= {16'd22400, 16'd23915};
                15'd7852 : data_rom <= {16'd22402, 16'd23913};
                15'd7853 : data_rom <= {16'd22405, 16'd23911};
                15'd7854 : data_rom <= {16'd22407, 16'd23909};
                15'd7855 : data_rom <= {16'd22409, 16'd23906};
                15'd7856 : data_rom <= {16'd22412, 16'd23904};
                15'd7857 : data_rom <= {16'd22414, 16'd23902};
                15'd7858 : data_rom <= {16'd22416, 16'd23900};
                15'd7859 : data_rom <= {16'd22419, 16'd23898};
                15'd7860 : data_rom <= {16'd22421, 16'd23896};
                15'd7861 : data_rom <= {16'd22423, 16'd23893};
                15'd7862 : data_rom <= {16'd22425, 16'd23891};
                15'd7863 : data_rom <= {16'd22428, 16'd23889};
                15'd7864 : data_rom <= {16'd22430, 16'd23887};
                15'd7865 : data_rom <= {16'd22432, 16'd23885};
                15'd7866 : data_rom <= {16'd22435, 16'd23883};
                15'd7867 : data_rom <= {16'd22437, 16'd23881};
                15'd7868 : data_rom <= {16'd22439, 16'd23878};
                15'd7869 : data_rom <= {16'd22441, 16'd23876};
                15'd7870 : data_rom <= {16'd22444, 16'd23874};
                15'd7871 : data_rom <= {16'd22446, 16'd23872};
                15'd7872 : data_rom <= {16'd22448, 16'd23870};
                15'd7873 : data_rom <= {16'd22451, 16'd23868};
                15'd7874 : data_rom <= {16'd22453, 16'd23866};
                15'd7875 : data_rom <= {16'd22455, 16'd23863};
                15'd7876 : data_rom <= {16'd22457, 16'd23861};
                15'd7877 : data_rom <= {16'd22460, 16'd23859};
                15'd7878 : data_rom <= {16'd22462, 16'd23857};
                15'd7879 : data_rom <= {16'd22464, 16'd23855};
                15'd7880 : data_rom <= {16'd22467, 16'd23853};
                15'd7881 : data_rom <= {16'd22469, 16'd23850};
                15'd7882 : data_rom <= {16'd22471, 16'd23848};
                15'd7883 : data_rom <= {16'd22473, 16'd23846};
                15'd7884 : data_rom <= {16'd22476, 16'd23844};
                15'd7885 : data_rom <= {16'd22478, 16'd23842};
                15'd7886 : data_rom <= {16'd22480, 16'd23840};
                15'd7887 : data_rom <= {16'd22483, 16'd23838};
                15'd7888 : data_rom <= {16'd22485, 16'd23835};
                15'd7889 : data_rom <= {16'd22487, 16'd23833};
                15'd7890 : data_rom <= {16'd22489, 16'd23831};
                15'd7891 : data_rom <= {16'd22492, 16'd23829};
                15'd7892 : data_rom <= {16'd22494, 16'd23827};
                15'd7893 : data_rom <= {16'd22496, 16'd23825};
                15'd7894 : data_rom <= {16'd22499, 16'd23822};
                15'd7895 : data_rom <= {16'd22501, 16'd23820};
                15'd7896 : data_rom <= {16'd22503, 16'd23818};
                15'd7897 : data_rom <= {16'd22505, 16'd23816};
                15'd7898 : data_rom <= {16'd22508, 16'd23814};
                15'd7899 : data_rom <= {16'd22510, 16'd23812};
                15'd7900 : data_rom <= {16'd22512, 16'd23809};
                15'd7901 : data_rom <= {16'd22515, 16'd23807};
                15'd7902 : data_rom <= {16'd22517, 16'd23805};
                15'd7903 : data_rom <= {16'd22519, 16'd23803};
                15'd7904 : data_rom <= {16'd22521, 16'd23801};
                15'd7905 : data_rom <= {16'd22524, 16'd23799};
                15'd7906 : data_rom <= {16'd22526, 16'd23797};
                15'd7907 : data_rom <= {16'd22528, 16'd23794};
                15'd7908 : data_rom <= {16'd22531, 16'd23792};
                15'd7909 : data_rom <= {16'd22533, 16'd23790};
                15'd7910 : data_rom <= {16'd22535, 16'd23788};
                15'd7911 : data_rom <= {16'd22537, 16'd23786};
                15'd7912 : data_rom <= {16'd22540, 16'd23784};
                15'd7913 : data_rom <= {16'd22542, 16'd23781};
                15'd7914 : data_rom <= {16'd22544, 16'd23779};
                15'd7915 : data_rom <= {16'd22547, 16'd23777};
                15'd7916 : data_rom <= {16'd22549, 16'd23775};
                15'd7917 : data_rom <= {16'd22551, 16'd23773};
                15'd7918 : data_rom <= {16'd22553, 16'd23771};
                15'd7919 : data_rom <= {16'd22556, 16'd23768};
                15'd7920 : data_rom <= {16'd22558, 16'd23766};
                15'd7921 : data_rom <= {16'd22560, 16'd23764};
                15'd7922 : data_rom <= {16'd22562, 16'd23762};
                15'd7923 : data_rom <= {16'd22565, 16'd23760};
                15'd7924 : data_rom <= {16'd22567, 16'd23758};
                15'd7925 : data_rom <= {16'd22569, 16'd23755};
                15'd7926 : data_rom <= {16'd22572, 16'd23753};
                15'd7927 : data_rom <= {16'd22574, 16'd23751};
                15'd7928 : data_rom <= {16'd22576, 16'd23749};
                15'd7929 : data_rom <= {16'd22578, 16'd23747};
                15'd7930 : data_rom <= {16'd22581, 16'd23745};
                15'd7931 : data_rom <= {16'd22583, 16'd23742};
                15'd7932 : data_rom <= {16'd22585, 16'd23740};
                15'd7933 : data_rom <= {16'd22588, 16'd23738};
                15'd7934 : data_rom <= {16'd22590, 16'd23736};
                15'd7935 : data_rom <= {16'd22592, 16'd23734};
                15'd7936 : data_rom <= {16'd22594, 16'd23732};
                15'd7937 : data_rom <= {16'd22597, 16'd23729};
                15'd7938 : data_rom <= {16'd22599, 16'd23727};
                15'd7939 : data_rom <= {16'd22601, 16'd23725};
                15'd7940 : data_rom <= {16'd22603, 16'd23723};
                15'd7941 : data_rom <= {16'd22606, 16'd23721};
                15'd7942 : data_rom <= {16'd22608, 16'd23719};
                15'd7943 : data_rom <= {16'd22610, 16'd23716};
                15'd7944 : data_rom <= {16'd22613, 16'd23714};
                15'd7945 : data_rom <= {16'd22615, 16'd23712};
                15'd7946 : data_rom <= {16'd22617, 16'd23710};
                15'd7947 : data_rom <= {16'd22619, 16'd23708};
                15'd7948 : data_rom <= {16'd22622, 16'd23706};
                15'd7949 : data_rom <= {16'd22624, 16'd23703};
                15'd7950 : data_rom <= {16'd22626, 16'd23701};
                15'd7951 : data_rom <= {16'd22628, 16'd23699};
                15'd7952 : data_rom <= {16'd22631, 16'd23697};
                15'd7953 : data_rom <= {16'd22633, 16'd23695};
                15'd7954 : data_rom <= {16'd22635, 16'd23693};
                15'd7955 : data_rom <= {16'd22638, 16'd23690};
                15'd7956 : data_rom <= {16'd22640, 16'd23688};
                15'd7957 : data_rom <= {16'd22642, 16'd23686};
                15'd7958 : data_rom <= {16'd22644, 16'd23684};
                15'd7959 : data_rom <= {16'd22647, 16'd23682};
                15'd7960 : data_rom <= {16'd22649, 16'd23680};
                15'd7961 : data_rom <= {16'd22651, 16'd23677};
                15'd7962 : data_rom <= {16'd22653, 16'd23675};
                15'd7963 : data_rom <= {16'd22656, 16'd23673};
                15'd7964 : data_rom <= {16'd22658, 16'd23671};
                15'd7965 : data_rom <= {16'd22660, 16'd23669};
                15'd7966 : data_rom <= {16'd22663, 16'd23667};
                15'd7967 : data_rom <= {16'd22665, 16'd23664};
                15'd7968 : data_rom <= {16'd22667, 16'd23662};
                15'd7969 : data_rom <= {16'd22669, 16'd23660};
                15'd7970 : data_rom <= {16'd22672, 16'd23658};
                15'd7971 : data_rom <= {16'd22674, 16'd23656};
                15'd7972 : data_rom <= {16'd22676, 16'd23654};
                15'd7973 : data_rom <= {16'd22678, 16'd23651};
                15'd7974 : data_rom <= {16'd22681, 16'd23649};
                15'd7975 : data_rom <= {16'd22683, 16'd23647};
                15'd7976 : data_rom <= {16'd22685, 16'd23645};
                15'd7977 : data_rom <= {16'd22687, 16'd23643};
                15'd7978 : data_rom <= {16'd22690, 16'd23640};
                15'd7979 : data_rom <= {16'd22692, 16'd23638};
                15'd7980 : data_rom <= {16'd22694, 16'd23636};
                15'd7981 : data_rom <= {16'd22697, 16'd23634};
                15'd7982 : data_rom <= {16'd22699, 16'd23632};
                15'd7983 : data_rom <= {16'd22701, 16'd23630};
                15'd7984 : data_rom <= {16'd22703, 16'd23627};
                15'd7985 : data_rom <= {16'd22706, 16'd23625};
                15'd7986 : data_rom <= {16'd22708, 16'd23623};
                15'd7987 : data_rom <= {16'd22710, 16'd23621};
                15'd7988 : data_rom <= {16'd22712, 16'd23619};
                15'd7989 : data_rom <= {16'd22715, 16'd23617};
                15'd7990 : data_rom <= {16'd22717, 16'd23614};
                15'd7991 : data_rom <= {16'd22719, 16'd23612};
                15'd7992 : data_rom <= {16'd22721, 16'd23610};
                15'd7993 : data_rom <= {16'd22724, 16'd23608};
                15'd7994 : data_rom <= {16'd22726, 16'd23606};
                15'd7995 : data_rom <= {16'd22728, 16'd23603};
                15'd7996 : data_rom <= {16'd22730, 16'd23601};
                15'd7997 : data_rom <= {16'd22733, 16'd23599};
                15'd7998 : data_rom <= {16'd22735, 16'd23597};
                15'd7999 : data_rom <= {16'd22737, 16'd23595};
                15'd8000 : data_rom <= {16'd22740, 16'd23593};
                15'd8001 : data_rom <= {16'd22742, 16'd23590};
                15'd8002 : data_rom <= {16'd22744, 16'd23588};
                15'd8003 : data_rom <= {16'd22746, 16'd23586};
                15'd8004 : data_rom <= {16'd22749, 16'd23584};
                15'd8005 : data_rom <= {16'd22751, 16'd23582};
                15'd8006 : data_rom <= {16'd22753, 16'd23579};
                15'd8007 : data_rom <= {16'd22755, 16'd23577};
                15'd8008 : data_rom <= {16'd22758, 16'd23575};
                15'd8009 : data_rom <= {16'd22760, 16'd23573};
                15'd8010 : data_rom <= {16'd22762, 16'd23571};
                15'd8011 : data_rom <= {16'd22764, 16'd23569};
                15'd8012 : data_rom <= {16'd22767, 16'd23566};
                15'd8013 : data_rom <= {16'd22769, 16'd23564};
                15'd8014 : data_rom <= {16'd22771, 16'd23562};
                15'd8015 : data_rom <= {16'd22773, 16'd23560};
                15'd8016 : data_rom <= {16'd22776, 16'd23558};
                15'd8017 : data_rom <= {16'd22778, 16'd23555};
                15'd8018 : data_rom <= {16'd22780, 16'd23553};
                15'd8019 : data_rom <= {16'd22782, 16'd23551};
                15'd8020 : data_rom <= {16'd22785, 16'd23549};
                15'd8021 : data_rom <= {16'd22787, 16'd23547};
                15'd8022 : data_rom <= {16'd22789, 16'd23545};
                15'd8023 : data_rom <= {16'd22792, 16'd23542};
                15'd8024 : data_rom <= {16'd22794, 16'd23540};
                15'd8025 : data_rom <= {16'd22796, 16'd23538};
                15'd8026 : data_rom <= {16'd22798, 16'd23536};
                15'd8027 : data_rom <= {16'd22801, 16'd23534};
                15'd8028 : data_rom <= {16'd22803, 16'd23531};
                15'd8029 : data_rom <= {16'd22805, 16'd23529};
                15'd8030 : data_rom <= {16'd22807, 16'd23527};
                15'd8031 : data_rom <= {16'd22810, 16'd23525};
                15'd8032 : data_rom <= {16'd22812, 16'd23523};
                15'd8033 : data_rom <= {16'd22814, 16'd23520};
                15'd8034 : data_rom <= {16'd22816, 16'd23518};
                15'd8035 : data_rom <= {16'd22819, 16'd23516};
                15'd8036 : data_rom <= {16'd22821, 16'd23514};
                15'd8037 : data_rom <= {16'd22823, 16'd23512};
                15'd8038 : data_rom <= {16'd22825, 16'd23510};
                15'd8039 : data_rom <= {16'd22828, 16'd23507};
                15'd8040 : data_rom <= {16'd22830, 16'd23505};
                15'd8041 : data_rom <= {16'd22832, 16'd23503};
                15'd8042 : data_rom <= {16'd22834, 16'd23501};
                15'd8043 : data_rom <= {16'd22837, 16'd23499};
                15'd8044 : data_rom <= {16'd22839, 16'd23496};
                15'd8045 : data_rom <= {16'd22841, 16'd23494};
                15'd8046 : data_rom <= {16'd22843, 16'd23492};
                15'd8047 : data_rom <= {16'd22846, 16'd23490};
                15'd8048 : data_rom <= {16'd22848, 16'd23488};
                15'd8049 : data_rom <= {16'd22850, 16'd23485};
                15'd8050 : data_rom <= {16'd22852, 16'd23483};
                15'd8051 : data_rom <= {16'd22855, 16'd23481};
                15'd8052 : data_rom <= {16'd22857, 16'd23479};
                15'd8053 : data_rom <= {16'd22859, 16'd23477};
                15'd8054 : data_rom <= {16'd22861, 16'd23475};
                15'd8055 : data_rom <= {16'd22864, 16'd23472};
                15'd8056 : data_rom <= {16'd22866, 16'd23470};
                15'd8057 : data_rom <= {16'd22868, 16'd23468};
                15'd8058 : data_rom <= {16'd22870, 16'd23466};
                15'd8059 : data_rom <= {16'd22873, 16'd23464};
                15'd8060 : data_rom <= {16'd22875, 16'd23461};
                15'd8061 : data_rom <= {16'd22877, 16'd23459};
                15'd8062 : data_rom <= {16'd22879, 16'd23457};
                15'd8063 : data_rom <= {16'd22882, 16'd23455};
                15'd8064 : data_rom <= {16'd22884, 16'd23453};
                15'd8065 : data_rom <= {16'd22886, 16'd23450};
                15'd8066 : data_rom <= {16'd22888, 16'd23448};
                15'd8067 : data_rom <= {16'd22891, 16'd23446};
                15'd8068 : data_rom <= {16'd22893, 16'd23444};
                15'd8069 : data_rom <= {16'd22895, 16'd23442};
                15'd8070 : data_rom <= {16'd22897, 16'd23439};
                15'd8071 : data_rom <= {16'd22900, 16'd23437};
                15'd8072 : data_rom <= {16'd22902, 16'd23435};
                15'd8073 : data_rom <= {16'd22904, 16'd23433};
                15'd8074 : data_rom <= {16'd22906, 16'd23431};
                15'd8075 : data_rom <= {16'd22909, 16'd23428};
                15'd8076 : data_rom <= {16'd22911, 16'd23426};
                15'd8077 : data_rom <= {16'd22913, 16'd23424};
                15'd8078 : data_rom <= {16'd22915, 16'd23422};
                15'd8079 : data_rom <= {16'd22918, 16'd23420};
                15'd8080 : data_rom <= {16'd22920, 16'd23417};
                15'd8081 : data_rom <= {16'd22922, 16'd23415};
                15'd8082 : data_rom <= {16'd22924, 16'd23413};
                15'd8083 : data_rom <= {16'd22927, 16'd23411};
                15'd8084 : data_rom <= {16'd22929, 16'd23409};
                15'd8085 : data_rom <= {16'd22931, 16'd23406};
                15'd8086 : data_rom <= {16'd22933, 16'd23404};
                15'd8087 : data_rom <= {16'd22936, 16'd23402};
                15'd8088 : data_rom <= {16'd22938, 16'd23400};
                15'd8089 : data_rom <= {16'd22940, 16'd23398};
                15'd8090 : data_rom <= {16'd22942, 16'd23395};
                15'd8091 : data_rom <= {16'd22945, 16'd23393};
                15'd8092 : data_rom <= {16'd22947, 16'd23391};
                15'd8093 : data_rom <= {16'd22949, 16'd23389};
                15'd8094 : data_rom <= {16'd22951, 16'd23387};
                15'd8095 : data_rom <= {16'd22953, 16'd23384};
                15'd8096 : data_rom <= {16'd22956, 16'd23382};
                15'd8097 : data_rom <= {16'd22958, 16'd23380};
                15'd8098 : data_rom <= {16'd22960, 16'd23378};
                15'd8099 : data_rom <= {16'd22962, 16'd23376};
                15'd8100 : data_rom <= {16'd22965, 16'd23373};
                15'd8101 : data_rom <= {16'd22967, 16'd23371};
                15'd8102 : data_rom <= {16'd22969, 16'd23369};
                15'd8103 : data_rom <= {16'd22971, 16'd23367};
                15'd8104 : data_rom <= {16'd22974, 16'd23365};
                15'd8105 : data_rom <= {16'd22976, 16'd23362};
                15'd8106 : data_rom <= {16'd22978, 16'd23360};
                15'd8107 : data_rom <= {16'd22980, 16'd23358};
                15'd8108 : data_rom <= {16'd22983, 16'd23356};
                15'd8109 : data_rom <= {16'd22985, 16'd23354};
                15'd8110 : data_rom <= {16'd22987, 16'd23351};
                15'd8111 : data_rom <= {16'd22989, 16'd23349};
                15'd8112 : data_rom <= {16'd22992, 16'd23347};
                15'd8113 : data_rom <= {16'd22994, 16'd23345};
                15'd8114 : data_rom <= {16'd22996, 16'd23343};
                15'd8115 : data_rom <= {16'd22998, 16'd23340};
                15'd8116 : data_rom <= {16'd23001, 16'd23338};
                15'd8117 : data_rom <= {16'd23003, 16'd23336};
                15'd8118 : data_rom <= {16'd23005, 16'd23334};
                15'd8119 : data_rom <= {16'd23007, 16'd23332};
                15'd8120 : data_rom <= {16'd23009, 16'd23329};
                15'd8121 : data_rom <= {16'd23012, 16'd23327};
                15'd8122 : data_rom <= {16'd23014, 16'd23325};
                15'd8123 : data_rom <= {16'd23016, 16'd23323};
                15'd8124 : data_rom <= {16'd23018, 16'd23321};
                15'd8125 : data_rom <= {16'd23021, 16'd23318};
                15'd8126 : data_rom <= {16'd23023, 16'd23316};
                15'd8127 : data_rom <= {16'd23025, 16'd23314};
                15'd8128 : data_rom <= {16'd23027, 16'd23312};
                15'd8129 : data_rom <= {16'd23030, 16'd23310};
                15'd8130 : data_rom <= {16'd23032, 16'd23307};
                15'd8131 : data_rom <= {16'd23034, 16'd23305};
                15'd8132 : data_rom <= {16'd23036, 16'd23303};
                15'd8133 : data_rom <= {16'd23039, 16'd23301};
                15'd8134 : data_rom <= {16'd23041, 16'd23298};
                15'd8135 : data_rom <= {16'd23043, 16'd23296};
                15'd8136 : data_rom <= {16'd23045, 16'd23294};
                15'd8137 : data_rom <= {16'd23047, 16'd23292};
                15'd8138 : data_rom <= {16'd23050, 16'd23290};
                15'd8139 : data_rom <= {16'd23052, 16'd23287};
                15'd8140 : data_rom <= {16'd23054, 16'd23285};
                15'd8141 : data_rom <= {16'd23056, 16'd23283};
                15'd8142 : data_rom <= {16'd23059, 16'd23281};
                15'd8143 : data_rom <= {16'd23061, 16'd23279};
                15'd8144 : data_rom <= {16'd23063, 16'd23276};
                15'd8145 : data_rom <= {16'd23065, 16'd23274};
                15'd8146 : data_rom <= {16'd23068, 16'd23272};
                15'd8147 : data_rom <= {16'd23070, 16'd23270};
                15'd8148 : data_rom <= {16'd23072, 16'd23268};
                15'd8149 : data_rom <= {16'd23074, 16'd23265};
                15'd8150 : data_rom <= {16'd23076, 16'd23263};
                15'd8151 : data_rom <= {16'd23079, 16'd23261};
                15'd8152 : data_rom <= {16'd23081, 16'd23259};
                15'd8153 : data_rom <= {16'd23083, 16'd23256};
                15'd8154 : data_rom <= {16'd23085, 16'd23254};
                15'd8155 : data_rom <= {16'd23088, 16'd23252};
                15'd8156 : data_rom <= {16'd23090, 16'd23250};
                15'd8157 : data_rom <= {16'd23092, 16'd23248};
                15'd8158 : data_rom <= {16'd23094, 16'd23245};
                15'd8159 : data_rom <= {16'd23097, 16'd23243};
                15'd8160 : data_rom <= {16'd23099, 16'd23241};
                15'd8161 : data_rom <= {16'd23101, 16'd23239};
                15'd8162 : data_rom <= {16'd23103, 16'd23237};
                15'd8163 : data_rom <= {16'd23105, 16'd23234};
                15'd8164 : data_rom <= {16'd23108, 16'd23232};
                15'd8165 : data_rom <= {16'd23110, 16'd23230};
                15'd8166 : data_rom <= {16'd23112, 16'd23228};
                15'd8167 : data_rom <= {16'd23114, 16'd23225};
                15'd8168 : data_rom <= {16'd23117, 16'd23223};
                15'd8169 : data_rom <= {16'd23119, 16'd23221};
                15'd8170 : data_rom <= {16'd23121, 16'd23219};
                15'd8171 : data_rom <= {16'd23123, 16'd23217};
                15'd8172 : data_rom <= {16'd23125, 16'd23214};
                15'd8173 : data_rom <= {16'd23128, 16'd23212};
                15'd8174 : data_rom <= {16'd23130, 16'd23210};
                15'd8175 : data_rom <= {16'd23132, 16'd23208};
                15'd8176 : data_rom <= {16'd23134, 16'd23206};
                15'd8177 : data_rom <= {16'd23137, 16'd23203};
                15'd8178 : data_rom <= {16'd23139, 16'd23201};
                15'd8179 : data_rom <= {16'd23141, 16'd23199};
                15'd8180 : data_rom <= {16'd23143, 16'd23197};
                15'd8181 : data_rom <= {16'd23146, 16'd23194};
                15'd8182 : data_rom <= {16'd23148, 16'd23192};
                15'd8183 : data_rom <= {16'd23150, 16'd23190};
                15'd8184 : data_rom <= {16'd23152, 16'd23188};
                15'd8185 : data_rom <= {16'd23154, 16'd23186};
                15'd8186 : data_rom <= {16'd23157, 16'd23183};
                15'd8187 : data_rom <= {16'd23159, 16'd23181};
                15'd8188 : data_rom <= {16'd23161, 16'd23179};
                15'd8189 : data_rom <= {16'd23163, 16'd23177};
                15'd8190 : data_rom <= {16'd23166, 16'd23174};
                15'd8191 : data_rom <= {16'd23168, 16'd23172};
                15'd8192 : data_rom <= {16'd23170, 16'd23170};
				15'd8193 : data_rom <= {16'd23172, 16'd23168};
                15'd8194 : data_rom <= {16'd23174, 16'd23166};
                15'd8195 : data_rom <= {16'd23177, 16'd23163};
                15'd8196 : data_rom <= {16'd23179, 16'd23161};
                15'd8197 : data_rom <= {16'd23181, 16'd23159};
                15'd8198 : data_rom <= {16'd23183, 16'd23157};
                15'd8199 : data_rom <= {16'd23186, 16'd23154};
                15'd8200 : data_rom <= {16'd23188, 16'd23152};
                15'd8201 : data_rom <= {16'd23190, 16'd23150};
                15'd8202 : data_rom <= {16'd23192, 16'd23148};
                15'd8203 : data_rom <= {16'd23194, 16'd23146};
                15'd8204 : data_rom <= {16'd23197, 16'd23143};
                15'd8205 : data_rom <= {16'd23199, 16'd23141};
                15'd8206 : data_rom <= {16'd23201, 16'd23139};
                15'd8207 : data_rom <= {16'd23203, 16'd23137};
                15'd8208 : data_rom <= {16'd23205, 16'd23134};
                15'd8209 : data_rom <= {16'd23208, 16'd23132};
                15'd8210 : data_rom <= {16'd23210, 16'd23130};
                15'd8211 : data_rom <= {16'd23212, 16'd23128};
                15'd8212 : data_rom <= {16'd23214, 16'd23126};
                15'd8213 : data_rom <= {16'd23217, 16'd23123};
                15'd8214 : data_rom <= {16'd23219, 16'd23121};
                15'd8215 : data_rom <= {16'd23221, 16'd23119};
                15'd8216 : data_rom <= {16'd23223, 16'd23117};
                15'd8217 : data_rom <= {16'd23225, 16'd23114};
                15'd8218 : data_rom <= {16'd23228, 16'd23112};
                15'd8219 : data_rom <= {16'd23230, 16'd23110};
                15'd8220 : data_rom <= {16'd23232, 16'd23108};
                15'd8221 : data_rom <= {16'd23234, 16'd23105};
                15'd8222 : data_rom <= {16'd23237, 16'd23103};
                15'd8223 : data_rom <= {16'd23239, 16'd23101};
                15'd8224 : data_rom <= {16'd23241, 16'd23099};
                15'd8225 : data_rom <= {16'd23243, 16'd23097};
                15'd8226 : data_rom <= {16'd23245, 16'd23094};
                15'd8227 : data_rom <= {16'd23248, 16'd23092};
                15'd8228 : data_rom <= {16'd23250, 16'd23090};
                15'd8229 : data_rom <= {16'd23252, 16'd23088};
                15'd8230 : data_rom <= {16'd23254, 16'd23085};
                15'd8231 : data_rom <= {16'd23256, 16'd23083};
                15'd8232 : data_rom <= {16'd23259, 16'd23081};
                15'd8233 : data_rom <= {16'd23261, 16'd23079};
                15'd8234 : data_rom <= {16'd23263, 16'd23077};
                15'd8235 : data_rom <= {16'd23265, 16'd23074};
                15'd8236 : data_rom <= {16'd23267, 16'd23072};
                15'd8237 : data_rom <= {16'd23270, 16'd23070};
                15'd8238 : data_rom <= {16'd23272, 16'd23068};
                15'd8239 : data_rom <= {16'd23274, 16'd23065};
                15'd8240 : data_rom <= {16'd23276, 16'd23063};
                15'd8241 : data_rom <= {16'd23279, 16'd23061};
                15'd8242 : data_rom <= {16'd23281, 16'd23059};
                15'd8243 : data_rom <= {16'd23283, 16'd23056};
                15'd8244 : data_rom <= {16'd23285, 16'd23054};
                15'd8245 : data_rom <= {16'd23287, 16'd23052};
                15'd8246 : data_rom <= {16'd23290, 16'd23050};
                15'd8247 : data_rom <= {16'd23292, 16'd23047};
                15'd8248 : data_rom <= {16'd23294, 16'd23045};
                15'd8249 : data_rom <= {16'd23296, 16'd23043};
                15'd8250 : data_rom <= {16'd23298, 16'd23041};
                15'd8251 : data_rom <= {16'd23301, 16'd23039};
                15'd8252 : data_rom <= {16'd23303, 16'd23036};
                15'd8253 : data_rom <= {16'd23305, 16'd23034};
                15'd8254 : data_rom <= {16'd23307, 16'd23032};
                15'd8255 : data_rom <= {16'd23309, 16'd23030};
                15'd8256 : data_rom <= {16'd23312, 16'd23027};
                15'd8257 : data_rom <= {16'd23314, 16'd23025};
                15'd8258 : data_rom <= {16'd23316, 16'd23023};
                15'd8259 : data_rom <= {16'd23318, 16'd23021};
                15'd8260 : data_rom <= {16'd23321, 16'd23018};
                15'd8261 : data_rom <= {16'd23323, 16'd23016};
                15'd8262 : data_rom <= {16'd23325, 16'd23014};
                15'd8263 : data_rom <= {16'd23327, 16'd23012};
                15'd8264 : data_rom <= {16'd23329, 16'd23009};
                15'd8265 : data_rom <= {16'd23332, 16'd23007};
                15'd8266 : data_rom <= {16'd23334, 16'd23005};
                15'd8267 : data_rom <= {16'd23336, 16'd23003};
                15'd8268 : data_rom <= {16'd23338, 16'd23001};
                15'd8269 : data_rom <= {16'd23340, 16'd22998};
                15'd8270 : data_rom <= {16'd23343, 16'd22996};
                15'd8271 : data_rom <= {16'd23345, 16'd22994};
                15'd8272 : data_rom <= {16'd23347, 16'd22992};
                15'd8273 : data_rom <= {16'd23349, 16'd22989};
                15'd8274 : data_rom <= {16'd23351, 16'd22987};
                15'd8275 : data_rom <= {16'd23354, 16'd22985};
                15'd8276 : data_rom <= {16'd23356, 16'd22983};
                15'd8277 : data_rom <= {16'd23358, 16'd22980};
                15'd8278 : data_rom <= {16'd23360, 16'd22978};
                15'd8279 : data_rom <= {16'd23362, 16'd22976};
                15'd8280 : data_rom <= {16'd23365, 16'd22974};
                15'd8281 : data_rom <= {16'd23367, 16'd22971};
                15'd8282 : data_rom <= {16'd23369, 16'd22969};
                15'd8283 : data_rom <= {16'd23371, 16'd22967};
                15'd8284 : data_rom <= {16'd23373, 16'd22965};
                15'd8285 : data_rom <= {16'd23376, 16'd22962};
                15'd8286 : data_rom <= {16'd23378, 16'd22960};
                15'd8287 : data_rom <= {16'd23380, 16'd22958};
                15'd8288 : data_rom <= {16'd23382, 16'd22956};
                15'd8289 : data_rom <= {16'd23384, 16'd22954};
                15'd8290 : data_rom <= {16'd23387, 16'd22951};
                15'd8291 : data_rom <= {16'd23389, 16'd22949};
                15'd8292 : data_rom <= {16'd23391, 16'd22947};
                15'd8293 : data_rom <= {16'd23393, 16'd22945};
                15'd8294 : data_rom <= {16'd23395, 16'd22942};
                15'd8295 : data_rom <= {16'd23398, 16'd22940};
                15'd8296 : data_rom <= {16'd23400, 16'd22938};
                15'd8297 : data_rom <= {16'd23402, 16'd22936};
                15'd8298 : data_rom <= {16'd23404, 16'd22933};
                15'd8299 : data_rom <= {16'd23406, 16'd22931};
                15'd8300 : data_rom <= {16'd23409, 16'd22929};
                15'd8301 : data_rom <= {16'd23411, 16'd22927};
                15'd8302 : data_rom <= {16'd23413, 16'd22924};
                15'd8303 : data_rom <= {16'd23415, 16'd22922};
                15'd8304 : data_rom <= {16'd23417, 16'd22920};
                15'd8305 : data_rom <= {16'd23420, 16'd22918};
                15'd8306 : data_rom <= {16'd23422, 16'd22915};
                15'd8307 : data_rom <= {16'd23424, 16'd22913};
                15'd8308 : data_rom <= {16'd23426, 16'd22911};
                15'd8309 : data_rom <= {16'd23428, 16'd22909};
                15'd8310 : data_rom <= {16'd23431, 16'd22906};
                15'd8311 : data_rom <= {16'd23433, 16'd22904};
                15'd8312 : data_rom <= {16'd23435, 16'd22902};
                15'd8313 : data_rom <= {16'd23437, 16'd22900};
                15'd8314 : data_rom <= {16'd23439, 16'd22897};
                15'd8315 : data_rom <= {16'd23442, 16'd22895};
                15'd8316 : data_rom <= {16'd23444, 16'd22893};
                15'd8317 : data_rom <= {16'd23446, 16'd22891};
                15'd8318 : data_rom <= {16'd23448, 16'd22888};
                15'd8319 : data_rom <= {16'd23450, 16'd22886};
                15'd8320 : data_rom <= {16'd23453, 16'd22884};
                15'd8321 : data_rom <= {16'd23455, 16'd22882};
                15'd8322 : data_rom <= {16'd23457, 16'd22879};
                15'd8323 : data_rom <= {16'd23459, 16'd22877};
                15'd8324 : data_rom <= {16'd23461, 16'd22875};
                15'd8325 : data_rom <= {16'd23464, 16'd22873};
                15'd8326 : data_rom <= {16'd23466, 16'd22870};
                15'd8327 : data_rom <= {16'd23468, 16'd22868};
                15'd8328 : data_rom <= {16'd23470, 16'd22866};
                15'd8329 : data_rom <= {16'd23472, 16'd22864};
                15'd8330 : data_rom <= {16'd23474, 16'd22861};
                15'd8331 : data_rom <= {16'd23477, 16'd22859};
                15'd8332 : data_rom <= {16'd23479, 16'd22857};
                15'd8333 : data_rom <= {16'd23481, 16'd22855};
                15'd8334 : data_rom <= {16'd23483, 16'd22852};
                15'd8335 : data_rom <= {16'd23485, 16'd22850};
                15'd8336 : data_rom <= {16'd23488, 16'd22848};
                15'd8337 : data_rom <= {16'd23490, 16'd22846};
                15'd8338 : data_rom <= {16'd23492, 16'd22843};
                15'd8339 : data_rom <= {16'd23494, 16'd22841};
                15'd8340 : data_rom <= {16'd23496, 16'd22839};
                15'd8341 : data_rom <= {16'd23499, 16'd22837};
                15'd8342 : data_rom <= {16'd23501, 16'd22834};
                15'd8343 : data_rom <= {16'd23503, 16'd22832};
                15'd8344 : data_rom <= {16'd23505, 16'd22830};
                15'd8345 : data_rom <= {16'd23507, 16'd22828};
                15'd8346 : data_rom <= {16'd23510, 16'd22825};
                15'd8347 : data_rom <= {16'd23512, 16'd22823};
                15'd8348 : data_rom <= {16'd23514, 16'd22821};
                15'd8349 : data_rom <= {16'd23516, 16'd22819};
                15'd8350 : data_rom <= {16'd23518, 16'd22816};
                15'd8351 : data_rom <= {16'd23520, 16'd22814};
                15'd8352 : data_rom <= {16'd23523, 16'd22812};
                15'd8353 : data_rom <= {16'd23525, 16'd22810};
                15'd8354 : data_rom <= {16'd23527, 16'd22807};
                15'd8355 : data_rom <= {16'd23529, 16'd22805};
                15'd8356 : data_rom <= {16'd23531, 16'd22803};
                15'd8357 : data_rom <= {16'd23534, 16'd22801};
                15'd8358 : data_rom <= {16'd23536, 16'd22798};
                15'd8359 : data_rom <= {16'd23538, 16'd22796};
                15'd8360 : data_rom <= {16'd23540, 16'd22794};
                15'd8361 : data_rom <= {16'd23542, 16'd22792};
                15'd8362 : data_rom <= {16'd23545, 16'd22789};
                15'd8363 : data_rom <= {16'd23547, 16'd22787};
                15'd8364 : data_rom <= {16'd23549, 16'd22785};
                15'd8365 : data_rom <= {16'd23551, 16'd22783};
                15'd8366 : data_rom <= {16'd23553, 16'd22780};
                15'd8367 : data_rom <= {16'd23555, 16'd22778};
                15'd8368 : data_rom <= {16'd23558, 16'd22776};
                15'd8369 : data_rom <= {16'd23560, 16'd22773};
                15'd8370 : data_rom <= {16'd23562, 16'd22771};
                15'd8371 : data_rom <= {16'd23564, 16'd22769};
                15'd8372 : data_rom <= {16'd23566, 16'd22767};
                15'd8373 : data_rom <= {16'd23569, 16'd22764};
                15'd8374 : data_rom <= {16'd23571, 16'd22762};
                15'd8375 : data_rom <= {16'd23573, 16'd22760};
                15'd8376 : data_rom <= {16'd23575, 16'd22758};
                15'd8377 : data_rom <= {16'd23577, 16'd22755};
                15'd8378 : data_rom <= {16'd23579, 16'd22753};
                15'd8379 : data_rom <= {16'd23582, 16'd22751};
                15'd8380 : data_rom <= {16'd23584, 16'd22749};
                15'd8381 : data_rom <= {16'd23586, 16'd22746};
                15'd8382 : data_rom <= {16'd23588, 16'd22744};
                15'd8383 : data_rom <= {16'd23590, 16'd22742};
                15'd8384 : data_rom <= {16'd23593, 16'd22740};
                15'd8385 : data_rom <= {16'd23595, 16'd22737};
                15'd8386 : data_rom <= {16'd23597, 16'd22735};
                15'd8387 : data_rom <= {16'd23599, 16'd22733};
                15'd8388 : data_rom <= {16'd23601, 16'd22731};
                15'd8389 : data_rom <= {16'd23603, 16'd22728};
                15'd8390 : data_rom <= {16'd23606, 16'd22726};
                15'd8391 : data_rom <= {16'd23608, 16'd22724};
                15'd8392 : data_rom <= {16'd23610, 16'd22721};
                15'd8393 : data_rom <= {16'd23612, 16'd22719};
                15'd8394 : data_rom <= {16'd23614, 16'd22717};
                15'd8395 : data_rom <= {16'd23616, 16'd22715};
                15'd8396 : data_rom <= {16'd23619, 16'd22712};
                15'd8397 : data_rom <= {16'd23621, 16'd22710};
                15'd8398 : data_rom <= {16'd23623, 16'd22708};
                15'd8399 : data_rom <= {16'd23625, 16'd22706};
                15'd8400 : data_rom <= {16'd23627, 16'd22703};
                15'd8401 : data_rom <= {16'd23630, 16'd22701};
                15'd8402 : data_rom <= {16'd23632, 16'd22699};
                15'd8403 : data_rom <= {16'd23634, 16'd22697};
                15'd8404 : data_rom <= {16'd23636, 16'd22694};
                15'd8405 : data_rom <= {16'd23638, 16'd22692};
                15'd8406 : data_rom <= {16'd23640, 16'd22690};
                15'd8407 : data_rom <= {16'd23643, 16'd22687};
                15'd8408 : data_rom <= {16'd23645, 16'd22685};
                15'd8409 : data_rom <= {16'd23647, 16'd22683};
                15'd8410 : data_rom <= {16'd23649, 16'd22681};
                15'd8411 : data_rom <= {16'd23651, 16'd22678};
                15'd8412 : data_rom <= {16'd23653, 16'd22676};
                15'd8413 : data_rom <= {16'd23656, 16'd22674};
                15'd8414 : data_rom <= {16'd23658, 16'd22672};
                15'd8415 : data_rom <= {16'd23660, 16'd22669};
                15'd8416 : data_rom <= {16'd23662, 16'd22667};
                15'd8417 : data_rom <= {16'd23664, 16'd22665};
                15'd8418 : data_rom <= {16'd23667, 16'd22663};
                15'd8419 : data_rom <= {16'd23669, 16'd22660};
                15'd8420 : data_rom <= {16'd23671, 16'd22658};
                15'd8421 : data_rom <= {16'd23673, 16'd22656};
                15'd8422 : data_rom <= {16'd23675, 16'd22653};
                15'd8423 : data_rom <= {16'd23677, 16'd22651};
                15'd8424 : data_rom <= {16'd23680, 16'd22649};
                15'd8425 : data_rom <= {16'd23682, 16'd22647};
                15'd8426 : data_rom <= {16'd23684, 16'd22644};
                15'd8427 : data_rom <= {16'd23686, 16'd22642};
                15'd8428 : data_rom <= {16'd23688, 16'd22640};
                15'd8429 : data_rom <= {16'd23690, 16'd22638};
                15'd8430 : data_rom <= {16'd23693, 16'd22635};
                15'd8431 : data_rom <= {16'd23695, 16'd22633};
                15'd8432 : data_rom <= {16'd23697, 16'd22631};
                15'd8433 : data_rom <= {16'd23699, 16'd22628};
                15'd8434 : data_rom <= {16'd23701, 16'd22626};
                15'd8435 : data_rom <= {16'd23703, 16'd22624};
                15'd8436 : data_rom <= {16'd23706, 16'd22622};
                15'd8437 : data_rom <= {16'd23708, 16'd22619};
                15'd8438 : data_rom <= {16'd23710, 16'd22617};
                15'd8439 : data_rom <= {16'd23712, 16'd22615};
                15'd8440 : data_rom <= {16'd23714, 16'd22613};
                15'd8441 : data_rom <= {16'd23716, 16'd22610};
                15'd8442 : data_rom <= {16'd23719, 16'd22608};
                15'd8443 : data_rom <= {16'd23721, 16'd22606};
                15'd8444 : data_rom <= {16'd23723, 16'd22603};
                15'd8445 : data_rom <= {16'd23725, 16'd22601};
                15'd8446 : data_rom <= {16'd23727, 16'd22599};
                15'd8447 : data_rom <= {16'd23729, 16'd22597};
                15'd8448 : data_rom <= {16'd23732, 16'd22594};
                15'd8449 : data_rom <= {16'd23734, 16'd22592};
                15'd8450 : data_rom <= {16'd23736, 16'd22590};
                15'd8451 : data_rom <= {16'd23738, 16'd22588};
                15'd8452 : data_rom <= {16'd23740, 16'd22585};
                15'd8453 : data_rom <= {16'd23742, 16'd22583};
                15'd8454 : data_rom <= {16'd23745, 16'd22581};
                15'd8455 : data_rom <= {16'd23747, 16'd22578};
                15'd8456 : data_rom <= {16'd23749, 16'd22576};
                15'd8457 : data_rom <= {16'd23751, 16'd22574};
                15'd8458 : data_rom <= {16'd23753, 16'd22572};
                15'd8459 : data_rom <= {16'd23755, 16'd22569};
                15'd8460 : data_rom <= {16'd23758, 16'd22567};
                15'd8461 : data_rom <= {16'd23760, 16'd22565};
                15'd8462 : data_rom <= {16'd23762, 16'd22563};
                15'd8463 : data_rom <= {16'd23764, 16'd22560};
                15'd8464 : data_rom <= {16'd23766, 16'd22558};
                15'd8465 : data_rom <= {16'd23768, 16'd22556};
                15'd8466 : data_rom <= {16'd23771, 16'd22553};
                15'd8467 : data_rom <= {16'd23773, 16'd22551};
                15'd8468 : data_rom <= {16'd23775, 16'd22549};
                15'd8469 : data_rom <= {16'd23777, 16'd22547};
                15'd8470 : data_rom <= {16'd23779, 16'd22544};
                15'd8471 : data_rom <= {16'd23781, 16'd22542};
                15'd8472 : data_rom <= {16'd23784, 16'd22540};
                15'd8473 : data_rom <= {16'd23786, 16'd22537};
                15'd8474 : data_rom <= {16'd23788, 16'd22535};
                15'd8475 : data_rom <= {16'd23790, 16'd22533};
                15'd8476 : data_rom <= {16'd23792, 16'd22531};
                15'd8477 : data_rom <= {16'd23794, 16'd22528};
                15'd8478 : data_rom <= {16'd23797, 16'd22526};
                15'd8479 : data_rom <= {16'd23799, 16'd22524};
                15'd8480 : data_rom <= {16'd23801, 16'd22521};
                15'd8481 : data_rom <= {16'd23803, 16'd22519};
                15'd8482 : data_rom <= {16'd23805, 16'd22517};
                15'd8483 : data_rom <= {16'd23807, 16'd22515};
                15'd8484 : data_rom <= {16'd23809, 16'd22512};
                15'd8485 : data_rom <= {16'd23812, 16'd22510};
                15'd8486 : data_rom <= {16'd23814, 16'd22508};
                15'd8487 : data_rom <= {16'd23816, 16'd22505};
                15'd8488 : data_rom <= {16'd23818, 16'd22503};
                15'd8489 : data_rom <= {16'd23820, 16'd22501};
                15'd8490 : data_rom <= {16'd23822, 16'd22499};
                15'd8491 : data_rom <= {16'd23825, 16'd22496};
                15'd8492 : data_rom <= {16'd23827, 16'd22494};
                15'd8493 : data_rom <= {16'd23829, 16'd22492};
                15'd8494 : data_rom <= {16'd23831, 16'd22490};
                15'd8495 : data_rom <= {16'd23833, 16'd22487};
                15'd8496 : data_rom <= {16'd23835, 16'd22485};
                15'd8497 : data_rom <= {16'd23837, 16'd22483};
                15'd8498 : data_rom <= {16'd23840, 16'd22480};
                15'd8499 : data_rom <= {16'd23842, 16'd22478};
                15'd8500 : data_rom <= {16'd23844, 16'd22476};
                15'd8501 : data_rom <= {16'd23846, 16'd22474};
                15'd8502 : data_rom <= {16'd23848, 16'd22471};
                15'd8503 : data_rom <= {16'd23850, 16'd22469};
                15'd8504 : data_rom <= {16'd23853, 16'd22467};
                15'd8505 : data_rom <= {16'd23855, 16'd22464};
                15'd8506 : data_rom <= {16'd23857, 16'd22462};
                15'd8507 : data_rom <= {16'd23859, 16'd22460};
                15'd8508 : data_rom <= {16'd23861, 16'd22457};
                15'd8509 : data_rom <= {16'd23863, 16'd22455};
                15'd8510 : data_rom <= {16'd23865, 16'd22453};
                15'd8511 : data_rom <= {16'd23868, 16'd22451};
                15'd8512 : data_rom <= {16'd23870, 16'd22448};
                15'd8513 : data_rom <= {16'd23872, 16'd22446};
                15'd8514 : data_rom <= {16'd23874, 16'd22444};
                15'd8515 : data_rom <= {16'd23876, 16'd22441};
                15'd8516 : data_rom <= {16'd23878, 16'd22439};
                15'd8517 : data_rom <= {16'd23881, 16'd22437};
                15'd8518 : data_rom <= {16'd23883, 16'd22435};
                15'd8519 : data_rom <= {16'd23885, 16'd22432};
                15'd8520 : data_rom <= {16'd23887, 16'd22430};
                15'd8521 : data_rom <= {16'd23889, 16'd22428};
                15'd8522 : data_rom <= {16'd23891, 16'd22425};
                15'd8523 : data_rom <= {16'd23893, 16'd22423};
                15'd8524 : data_rom <= {16'd23896, 16'd22421};
                15'd8525 : data_rom <= {16'd23898, 16'd22419};
                15'd8526 : data_rom <= {16'd23900, 16'd22416};
                15'd8527 : data_rom <= {16'd23902, 16'd22414};
                15'd8528 : data_rom <= {16'd23904, 16'd22412};
                15'd8529 : data_rom <= {16'd23906, 16'd22409};
                15'd8530 : data_rom <= {16'd23909, 16'd22407};
                15'd8531 : data_rom <= {16'd23911, 16'd22405};
                15'd8532 : data_rom <= {16'd23913, 16'd22403};
                15'd8533 : data_rom <= {16'd23915, 16'd22400};
                15'd8534 : data_rom <= {16'd23917, 16'd22398};
                15'd8535 : data_rom <= {16'd23919, 16'd22396};
                15'd8536 : data_rom <= {16'd23921, 16'd22393};
                15'd8537 : data_rom <= {16'd23924, 16'd22391};
                15'd8538 : data_rom <= {16'd23926, 16'd22389};
                15'd8539 : data_rom <= {16'd23928, 16'd22386};
                15'd8540 : data_rom <= {16'd23930, 16'd22384};
                15'd8541 : data_rom <= {16'd23932, 16'd22382};
                15'd8542 : data_rom <= {16'd23934, 16'd22380};
                15'd8543 : data_rom <= {16'd23936, 16'd22377};
                15'd8544 : data_rom <= {16'd23939, 16'd22375};
                15'd8545 : data_rom <= {16'd23941, 16'd22373};
                15'd8546 : data_rom <= {16'd23943, 16'd22370};
                15'd8547 : data_rom <= {16'd23945, 16'd22368};
                15'd8548 : data_rom <= {16'd23947, 16'd22366};
                15'd8549 : data_rom <= {16'd23949, 16'd22364};
                15'd8550 : data_rom <= {16'd23951, 16'd22361};
                15'd8551 : data_rom <= {16'd23954, 16'd22359};
                15'd8552 : data_rom <= {16'd23956, 16'd22357};
                15'd8553 : data_rom <= {16'd23958, 16'd22354};
                15'd8554 : data_rom <= {16'd23960, 16'd22352};
                15'd8555 : data_rom <= {16'd23962, 16'd22350};
                15'd8556 : data_rom <= {16'd23964, 16'd22347};
                15'd8557 : data_rom <= {16'd23966, 16'd22345};
                15'd8558 : data_rom <= {16'd23969, 16'd22343};
                15'd8559 : data_rom <= {16'd23971, 16'd22341};
                15'd8560 : data_rom <= {16'd23973, 16'd22338};
                15'd8561 : data_rom <= {16'd23975, 16'd22336};
                15'd8562 : data_rom <= {16'd23977, 16'd22334};
                15'd8563 : data_rom <= {16'd23979, 16'd22331};
                15'd8564 : data_rom <= {16'd23981, 16'd22329};
                15'd8565 : data_rom <= {16'd23984, 16'd22327};
                15'd8566 : data_rom <= {16'd23986, 16'd22324};
                15'd8567 : data_rom <= {16'd23988, 16'd22322};
                15'd8568 : data_rom <= {16'd23990, 16'd22320};
                15'd8569 : data_rom <= {16'd23992, 16'd22318};
                15'd8570 : data_rom <= {16'd23994, 16'd22315};
                15'd8571 : data_rom <= {16'd23996, 16'd22313};
                15'd8572 : data_rom <= {16'd23999, 16'd22311};
                15'd8573 : data_rom <= {16'd24001, 16'd22308};
                15'd8574 : data_rom <= {16'd24003, 16'd22306};
                15'd8575 : data_rom <= {16'd24005, 16'd22304};
                15'd8576 : data_rom <= {16'd24007, 16'd22301};
                15'd8577 : data_rom <= {16'd24009, 16'd22299};
                15'd8578 : data_rom <= {16'd24011, 16'd22297};
                15'd8579 : data_rom <= {16'd24014, 16'd22295};
                15'd8580 : data_rom <= {16'd24016, 16'd22292};
                15'd8581 : data_rom <= {16'd24018, 16'd22290};
                15'd8582 : data_rom <= {16'd24020, 16'd22288};
                15'd8583 : data_rom <= {16'd24022, 16'd22285};
                15'd8584 : data_rom <= {16'd24024, 16'd22283};
                15'd8585 : data_rom <= {16'd24026, 16'd22281};
                15'd8586 : data_rom <= {16'd24028, 16'd22278};
                15'd8587 : data_rom <= {16'd24031, 16'd22276};
                15'd8588 : data_rom <= {16'd24033, 16'd22274};
                15'd8589 : data_rom <= {16'd24035, 16'd22272};
                15'd8590 : data_rom <= {16'd24037, 16'd22269};
                15'd8591 : data_rom <= {16'd24039, 16'd22267};
                15'd8592 : data_rom <= {16'd24041, 16'd22265};
                15'd8593 : data_rom <= {16'd24043, 16'd22262};
                15'd8594 : data_rom <= {16'd24046, 16'd22260};
                15'd8595 : data_rom <= {16'd24048, 16'd22258};
                15'd8596 : data_rom <= {16'd24050, 16'd22255};
                15'd8597 : data_rom <= {16'd24052, 16'd22253};
                15'd8598 : data_rom <= {16'd24054, 16'd22251};
                15'd8599 : data_rom <= {16'd24056, 16'd22248};
                15'd8600 : data_rom <= {16'd24058, 16'd22246};
                15'd8601 : data_rom <= {16'd24060, 16'd22244};
                15'd8602 : data_rom <= {16'd24063, 16'd22242};
                15'd8603 : data_rom <= {16'd24065, 16'd22239};
                15'd8604 : data_rom <= {16'd24067, 16'd22237};
                15'd8605 : data_rom <= {16'd24069, 16'd22235};
                15'd8606 : data_rom <= {16'd24071, 16'd22232};
                15'd8607 : data_rom <= {16'd24073, 16'd22230};
                15'd8608 : data_rom <= {16'd24075, 16'd22228};
                15'd8609 : data_rom <= {16'd24078, 16'd22225};
                15'd8610 : data_rom <= {16'd24080, 16'd22223};
                15'd8611 : data_rom <= {16'd24082, 16'd22221};
                15'd8612 : data_rom <= {16'd24084, 16'd22218};
                15'd8613 : data_rom <= {16'd24086, 16'd22216};
                15'd8614 : data_rom <= {16'd24088, 16'd22214};
                15'd8615 : data_rom <= {16'd24090, 16'd22212};
                15'd8616 : data_rom <= {16'd24092, 16'd22209};
                15'd8617 : data_rom <= {16'd24095, 16'd22207};
                15'd8618 : data_rom <= {16'd24097, 16'd22205};
                15'd8619 : data_rom <= {16'd24099, 16'd22202};
                15'd8620 : data_rom <= {16'd24101, 16'd22200};
                15'd8621 : data_rom <= {16'd24103, 16'd22198};
                15'd8622 : data_rom <= {16'd24105, 16'd22195};
                15'd8623 : data_rom <= {16'd24107, 16'd22193};
                15'd8624 : data_rom <= {16'd24109, 16'd22191};
                15'd8625 : data_rom <= {16'd24112, 16'd22188};
                15'd8626 : data_rom <= {16'd24114, 16'd22186};
                15'd8627 : data_rom <= {16'd24116, 16'd22184};
                15'd8628 : data_rom <= {16'd24118, 16'd22181};
                15'd8629 : data_rom <= {16'd24120, 16'd22179};
                15'd8630 : data_rom <= {16'd24122, 16'd22177};
                15'd8631 : data_rom <= {16'd24124, 16'd22175};
                15'd8632 : data_rom <= {16'd24126, 16'd22172};
                15'd8633 : data_rom <= {16'd24129, 16'd22170};
                15'd8634 : data_rom <= {16'd24131, 16'd22168};
                15'd8635 : data_rom <= {16'd24133, 16'd22165};
                15'd8636 : data_rom <= {16'd24135, 16'd22163};
                15'd8637 : data_rom <= {16'd24137, 16'd22161};
                15'd8638 : data_rom <= {16'd24139, 16'd22158};
                15'd8639 : data_rom <= {16'd24141, 16'd22156};
                15'd8640 : data_rom <= {16'd24143, 16'd22154};
                15'd8641 : data_rom <= {16'd24146, 16'd22151};
                15'd8642 : data_rom <= {16'd24148, 16'd22149};
                15'd8643 : data_rom <= {16'd24150, 16'd22147};
                15'd8644 : data_rom <= {16'd24152, 16'd22144};
                15'd8645 : data_rom <= {16'd24154, 16'd22142};
                15'd8646 : data_rom <= {16'd24156, 16'd22140};
                15'd8647 : data_rom <= {16'd24158, 16'd22138};
                15'd8648 : data_rom <= {16'd24160, 16'd22135};
                15'd8649 : data_rom <= {16'd24163, 16'd22133};
                15'd8650 : data_rom <= {16'd24165, 16'd22131};
                15'd8651 : data_rom <= {16'd24167, 16'd22128};
                15'd8652 : data_rom <= {16'd24169, 16'd22126};
                15'd8653 : data_rom <= {16'd24171, 16'd22124};
                15'd8654 : data_rom <= {16'd24173, 16'd22121};
                15'd8655 : data_rom <= {16'd24175, 16'd22119};
                15'd8656 : data_rom <= {16'd24177, 16'd22117};
                15'd8657 : data_rom <= {16'd24180, 16'd22114};
                15'd8658 : data_rom <= {16'd24182, 16'd22112};
                15'd8659 : data_rom <= {16'd24184, 16'd22110};
                15'd8660 : data_rom <= {16'd24186, 16'd22107};
                15'd8661 : data_rom <= {16'd24188, 16'd22105};
                15'd8662 : data_rom <= {16'd24190, 16'd22103};
                15'd8663 : data_rom <= {16'd24192, 16'd22100};
                15'd8664 : data_rom <= {16'd24194, 16'd22098};
                15'd8665 : data_rom <= {16'd24197, 16'd22096};
                15'd8666 : data_rom <= {16'd24199, 16'd22093};
                15'd8667 : data_rom <= {16'd24201, 16'd22091};
                15'd8668 : data_rom <= {16'd24203, 16'd22089};
                15'd8669 : data_rom <= {16'd24205, 16'd22087};
                15'd8670 : data_rom <= {16'd24207, 16'd22084};
                15'd8671 : data_rom <= {16'd24209, 16'd22082};
                15'd8672 : data_rom <= {16'd24211, 16'd22080};
                15'd8673 : data_rom <= {16'd24213, 16'd22077};
                15'd8674 : data_rom <= {16'd24216, 16'd22075};
                15'd8675 : data_rom <= {16'd24218, 16'd22073};
                15'd8676 : data_rom <= {16'd24220, 16'd22070};
                15'd8677 : data_rom <= {16'd24222, 16'd22068};
                15'd8678 : data_rom <= {16'd24224, 16'd22066};
                15'd8679 : data_rom <= {16'd24226, 16'd22063};
                15'd8680 : data_rom <= {16'd24228, 16'd22061};
                15'd8681 : data_rom <= {16'd24230, 16'd22059};
                15'd8682 : data_rom <= {16'd24233, 16'd22056};
                15'd8683 : data_rom <= {16'd24235, 16'd22054};
                15'd8684 : data_rom <= {16'd24237, 16'd22052};
                15'd8685 : data_rom <= {16'd24239, 16'd22049};
                15'd8686 : data_rom <= {16'd24241, 16'd22047};
                15'd8687 : data_rom <= {16'd24243, 16'd22045};
                15'd8688 : data_rom <= {16'd24245, 16'd22042};
                15'd8689 : data_rom <= {16'd24247, 16'd22040};
                15'd8690 : data_rom <= {16'd24249, 16'd22038};
                15'd8691 : data_rom <= {16'd24252, 16'd22035};
                15'd8692 : data_rom <= {16'd24254, 16'd22033};
                15'd8693 : data_rom <= {16'd24256, 16'd22031};
                15'd8694 : data_rom <= {16'd24258, 16'd22028};
                15'd8695 : data_rom <= {16'd24260, 16'd22026};
                15'd8696 : data_rom <= {16'd24262, 16'd22024};
                15'd8697 : data_rom <= {16'd24264, 16'd22021};
                15'd8698 : data_rom <= {16'd24266, 16'd22019};
                15'd8699 : data_rom <= {16'd24268, 16'd22017};
                15'd8700 : data_rom <= {16'd24271, 16'd22014};
                15'd8701 : data_rom <= {16'd24273, 16'd22012};
                15'd8702 : data_rom <= {16'd24275, 16'd22010};
                15'd8703 : data_rom <= {16'd24277, 16'd22007};
                15'd8704 : data_rom <= {16'd24279, 16'd22005};
                15'd8705 : data_rom <= {16'd24281, 16'd22003};
                15'd8706 : data_rom <= {16'd24283, 16'd22001};
                15'd8707 : data_rom <= {16'd24285, 16'd21998};
                15'd8708 : data_rom <= {16'd24287, 16'd21996};
                15'd8709 : data_rom <= {16'd24290, 16'd21994};
                15'd8710 : data_rom <= {16'd24292, 16'd21991};
                15'd8711 : data_rom <= {16'd24294, 16'd21989};
                15'd8712 : data_rom <= {16'd24296, 16'd21987};
                15'd8713 : data_rom <= {16'd24298, 16'd21984};
                15'd8714 : data_rom <= {16'd24300, 16'd21982};
                15'd8715 : data_rom <= {16'd24302, 16'd21980};
                15'd8716 : data_rom <= {16'd24304, 16'd21977};
                15'd8717 : data_rom <= {16'd24306, 16'd21975};
                15'd8718 : data_rom <= {16'd24308, 16'd21973};
                15'd8719 : data_rom <= {16'd24311, 16'd21970};
                15'd8720 : data_rom <= {16'd24313, 16'd21968};
                15'd8721 : data_rom <= {16'd24315, 16'd21966};
                15'd8722 : data_rom <= {16'd24317, 16'd21963};
                15'd8723 : data_rom <= {16'd24319, 16'd21961};
                15'd8724 : data_rom <= {16'd24321, 16'd21959};
                15'd8725 : data_rom <= {16'd24323, 16'd21956};
                15'd8726 : data_rom <= {16'd24325, 16'd21954};
                15'd8727 : data_rom <= {16'd24327, 16'd21952};
                15'd8728 : data_rom <= {16'd24330, 16'd21949};
                15'd8729 : data_rom <= {16'd24332, 16'd21947};
                15'd8730 : data_rom <= {16'd24334, 16'd21945};
                15'd8731 : data_rom <= {16'd24336, 16'd21942};
                15'd8732 : data_rom <= {16'd24338, 16'd21940};
                15'd8733 : data_rom <= {16'd24340, 16'd21938};
                15'd8734 : data_rom <= {16'd24342, 16'd21935};
                15'd8735 : data_rom <= {16'd24344, 16'd21933};
                15'd8736 : data_rom <= {16'd24346, 16'd21931};
                15'd8737 : data_rom <= {16'd24348, 16'd21928};
                15'd8738 : data_rom <= {16'd24351, 16'd21926};
                15'd8739 : data_rom <= {16'd24353, 16'd21924};
                15'd8740 : data_rom <= {16'd24355, 16'd21921};
                15'd8741 : data_rom <= {16'd24357, 16'd21919};
                15'd8742 : data_rom <= {16'd24359, 16'd21917};
                15'd8743 : data_rom <= {16'd24361, 16'd21914};
                15'd8744 : data_rom <= {16'd24363, 16'd21912};
                15'd8745 : data_rom <= {16'd24365, 16'd21910};
                15'd8746 : data_rom <= {16'd24367, 16'd21907};
                15'd8747 : data_rom <= {16'd24369, 16'd21905};
                15'd8748 : data_rom <= {16'd24372, 16'd21903};
                15'd8749 : data_rom <= {16'd24374, 16'd21900};
                15'd8750 : data_rom <= {16'd24376, 16'd21898};
                15'd8751 : data_rom <= {16'd24378, 16'd21896};
                15'd8752 : data_rom <= {16'd24380, 16'd21893};
                15'd8753 : data_rom <= {16'd24382, 16'd21891};
                15'd8754 : data_rom <= {16'd24384, 16'd21889};
                15'd8755 : data_rom <= {16'd24386, 16'd21886};
                15'd8756 : data_rom <= {16'd24388, 16'd21884};
                15'd8757 : data_rom <= {16'd24390, 16'd21882};
                15'd8758 : data_rom <= {16'd24393, 16'd21879};
                15'd8759 : data_rom <= {16'd24395, 16'd21877};
                15'd8760 : data_rom <= {16'd24397, 16'd21874};
                15'd8761 : data_rom <= {16'd24399, 16'd21872};
                15'd8762 : data_rom <= {16'd24401, 16'd21870};
                15'd8763 : data_rom <= {16'd24403, 16'd21867};
                15'd8764 : data_rom <= {16'd24405, 16'd21865};
                15'd8765 : data_rom <= {16'd24407, 16'd21863};
                15'd8766 : data_rom <= {16'd24409, 16'd21860};
                15'd8767 : data_rom <= {16'd24411, 16'd21858};
                15'd8768 : data_rom <= {16'd24414, 16'd21856};
                15'd8769 : data_rom <= {16'd24416, 16'd21853};
                15'd8770 : data_rom <= {16'd24418, 16'd21851};
                15'd8771 : data_rom <= {16'd24420, 16'd21849};
                15'd8772 : data_rom <= {16'd24422, 16'd21846};
                15'd8773 : data_rom <= {16'd24424, 16'd21844};
                15'd8774 : data_rom <= {16'd24426, 16'd21842};
                15'd8775 : data_rom <= {16'd24428, 16'd21839};
                15'd8776 : data_rom <= {16'd24430, 16'd21837};
                15'd8777 : data_rom <= {16'd24432, 16'd21835};
                15'd8778 : data_rom <= {16'd24434, 16'd21832};
                15'd8779 : data_rom <= {16'd24437, 16'd21830};
                15'd8780 : data_rom <= {16'd24439, 16'd21828};
                15'd8781 : data_rom <= {16'd24441, 16'd21825};
                15'd8782 : data_rom <= {16'd24443, 16'd21823};
                15'd8783 : data_rom <= {16'd24445, 16'd21821};
                15'd8784 : data_rom <= {16'd24447, 16'd21818};
                15'd8785 : data_rom <= {16'd24449, 16'd21816};
                15'd8786 : data_rom <= {16'd24451, 16'd21814};
                15'd8787 : data_rom <= {16'd24453, 16'd21811};
                15'd8788 : data_rom <= {16'd24455, 16'd21809};
                15'd8789 : data_rom <= {16'd24457, 16'd21807};
                15'd8790 : data_rom <= {16'd24460, 16'd21804};
                15'd8791 : data_rom <= {16'd24462, 16'd21802};
                15'd8792 : data_rom <= {16'd24464, 16'd21800};
                15'd8793 : data_rom <= {16'd24466, 16'd21797};
                15'd8794 : data_rom <= {16'd24468, 16'd21795};
                15'd8795 : data_rom <= {16'd24470, 16'd21793};
                15'd8796 : data_rom <= {16'd24472, 16'd21790};
                15'd8797 : data_rom <= {16'd24474, 16'd21788};
                15'd8798 : data_rom <= {16'd24476, 16'd21785};
                15'd8799 : data_rom <= {16'd24478, 16'd21783};
                15'd8800 : data_rom <= {16'd24480, 16'd21781};
                15'd8801 : data_rom <= {16'd24483, 16'd21778};
                15'd8802 : data_rom <= {16'd24485, 16'd21776};
                15'd8803 : data_rom <= {16'd24487, 16'd21774};
                15'd8804 : data_rom <= {16'd24489, 16'd21771};
                15'd8805 : data_rom <= {16'd24491, 16'd21769};
                15'd8806 : data_rom <= {16'd24493, 16'd21767};
                15'd8807 : data_rom <= {16'd24495, 16'd21764};
                15'd8808 : data_rom <= {16'd24497, 16'd21762};
                15'd8809 : data_rom <= {16'd24499, 16'd21760};
                15'd8810 : data_rom <= {16'd24501, 16'd21757};
                15'd8811 : data_rom <= {16'd24503, 16'd21755};
                15'd8812 : data_rom <= {16'd24506, 16'd21753};
                15'd8813 : data_rom <= {16'd24508, 16'd21750};
                15'd8814 : data_rom <= {16'd24510, 16'd21748};
                15'd8815 : data_rom <= {16'd24512, 16'd21746};
                15'd8816 : data_rom <= {16'd24514, 16'd21743};
                15'd8817 : data_rom <= {16'd24516, 16'd21741};
                15'd8818 : data_rom <= {16'd24518, 16'd21738};
                15'd8819 : data_rom <= {16'd24520, 16'd21736};
                15'd8820 : data_rom <= {16'd24522, 16'd21734};
                15'd8821 : data_rom <= {16'd24524, 16'd21731};
                15'd8822 : data_rom <= {16'd24526, 16'd21729};
                15'd8823 : data_rom <= {16'd24528, 16'd21727};
                15'd8824 : data_rom <= {16'd24531, 16'd21724};
                15'd8825 : data_rom <= {16'd24533, 16'd21722};
                15'd8826 : data_rom <= {16'd24535, 16'd21720};
                15'd8827 : data_rom <= {16'd24537, 16'd21717};
                15'd8828 : data_rom <= {16'd24539, 16'd21715};
                15'd8829 : data_rom <= {16'd24541, 16'd21713};
                15'd8830 : data_rom <= {16'd24543, 16'd21710};
                15'd8831 : data_rom <= {16'd24545, 16'd21708};
                15'd8832 : data_rom <= {16'd24547, 16'd21706};
                15'd8833 : data_rom <= {16'd24549, 16'd21703};
                15'd8834 : data_rom <= {16'd24551, 16'd21701};
                15'd8835 : data_rom <= {16'd24553, 16'd21698};
                15'd8836 : data_rom <= {16'd24556, 16'd21696};
                15'd8837 : data_rom <= {16'd24558, 16'd21694};
                15'd8838 : data_rom <= {16'd24560, 16'd21691};
                15'd8839 : data_rom <= {16'd24562, 16'd21689};
                15'd8840 : data_rom <= {16'd24564, 16'd21687};
                15'd8841 : data_rom <= {16'd24566, 16'd21684};
                15'd8842 : data_rom <= {16'd24568, 16'd21682};
                15'd8843 : data_rom <= {16'd24570, 16'd21680};
                15'd8844 : data_rom <= {16'd24572, 16'd21677};
                15'd8845 : data_rom <= {16'd24574, 16'd21675};
                15'd8846 : data_rom <= {16'd24576, 16'd21673};
                15'd8847 : data_rom <= {16'd24578, 16'd21670};
                15'd8848 : data_rom <= {16'd24580, 16'd21668};
                15'd8849 : data_rom <= {16'd24583, 16'd21666};
                15'd8850 : data_rom <= {16'd24585, 16'd21663};
                15'd8851 : data_rom <= {16'd24587, 16'd21661};
                15'd8852 : data_rom <= {16'd24589, 16'd21658};
                15'd8853 : data_rom <= {16'd24591, 16'd21656};
                15'd8854 : data_rom <= {16'd24593, 16'd21654};
                15'd8855 : data_rom <= {16'd24595, 16'd21651};
                15'd8856 : data_rom <= {16'd24597, 16'd21649};
                15'd8857 : data_rom <= {16'd24599, 16'd21647};
                15'd8858 : data_rom <= {16'd24601, 16'd21644};
                15'd8859 : data_rom <= {16'd24603, 16'd21642};
                15'd8860 : data_rom <= {16'd24605, 16'd21640};
                15'd8861 : data_rom <= {16'd24607, 16'd21637};
                15'd8862 : data_rom <= {16'd24610, 16'd21635};
                15'd8863 : data_rom <= {16'd24612, 16'd21633};
                15'd8864 : data_rom <= {16'd24614, 16'd21630};
                15'd8865 : data_rom <= {16'd24616, 16'd21628};
                15'd8866 : data_rom <= {16'd24618, 16'd21625};
                15'd8867 : data_rom <= {16'd24620, 16'd21623};
                15'd8868 : data_rom <= {16'd24622, 16'd21621};
                15'd8869 : data_rom <= {16'd24624, 16'd21618};
                15'd8870 : data_rom <= {16'd24626, 16'd21616};
                15'd8871 : data_rom <= {16'd24628, 16'd21614};
                15'd8872 : data_rom <= {16'd24630, 16'd21611};
                15'd8873 : data_rom <= {16'd24632, 16'd21609};
                15'd8874 : data_rom <= {16'd24634, 16'd21607};
                15'd8875 : data_rom <= {16'd24636, 16'd21604};
                15'd8876 : data_rom <= {16'd24639, 16'd21602};
                15'd8877 : data_rom <= {16'd24641, 16'd21599};
                15'd8878 : data_rom <= {16'd24643, 16'd21597};
                15'd8879 : data_rom <= {16'd24645, 16'd21595};
                15'd8880 : data_rom <= {16'd24647, 16'd21592};
                15'd8881 : data_rom <= {16'd24649, 16'd21590};
                15'd8882 : data_rom <= {16'd24651, 16'd21588};
                15'd8883 : data_rom <= {16'd24653, 16'd21585};
                15'd8884 : data_rom <= {16'd24655, 16'd21583};
                15'd8885 : data_rom <= {16'd24657, 16'd21581};
                15'd8886 : data_rom <= {16'd24659, 16'd21578};
                15'd8887 : data_rom <= {16'd24661, 16'd21576};
                15'd8888 : data_rom <= {16'd24663, 16'd21573};
                15'd8889 : data_rom <= {16'd24665, 16'd21571};
                15'd8890 : data_rom <= {16'd24668, 16'd21569};
                15'd8891 : data_rom <= {16'd24670, 16'd21566};
                15'd8892 : data_rom <= {16'd24672, 16'd21564};
                15'd8893 : data_rom <= {16'd24674, 16'd21562};
                15'd8894 : data_rom <= {16'd24676, 16'd21559};
                15'd8895 : data_rom <= {16'd24678, 16'd21557};
                15'd8896 : data_rom <= {16'd24680, 16'd21555};
                15'd8897 : data_rom <= {16'd24682, 16'd21552};
                15'd8898 : data_rom <= {16'd24684, 16'd21550};
                15'd8899 : data_rom <= {16'd24686, 16'd21547};
                15'd8900 : data_rom <= {16'd24688, 16'd21545};
                15'd8901 : data_rom <= {16'd24690, 16'd21543};
                15'd8902 : data_rom <= {16'd24692, 16'd21540};
                15'd8903 : data_rom <= {16'd24694, 16'd21538};
                15'd8904 : data_rom <= {16'd24696, 16'd21536};
                15'd8905 : data_rom <= {16'd24698, 16'd21533};
                15'd8906 : data_rom <= {16'd24701, 16'd21531};
                15'd8907 : data_rom <= {16'd24703, 16'd21528};
                15'd8908 : data_rom <= {16'd24705, 16'd21526};
                15'd8909 : data_rom <= {16'd24707, 16'd21524};
                15'd8910 : data_rom <= {16'd24709, 16'd21521};
                15'd8911 : data_rom <= {16'd24711, 16'd21519};
                15'd8912 : data_rom <= {16'd24713, 16'd21517};
                15'd8913 : data_rom <= {16'd24715, 16'd21514};
                15'd8914 : data_rom <= {16'd24717, 16'd21512};
                15'd8915 : data_rom <= {16'd24719, 16'd21510};
                15'd8916 : data_rom <= {16'd24721, 16'd21507};
                15'd8917 : data_rom <= {16'd24723, 16'd21505};
                15'd8918 : data_rom <= {16'd24725, 16'd21502};
                15'd8919 : data_rom <= {16'd24727, 16'd21500};
                15'd8920 : data_rom <= {16'd24729, 16'd21498};
                15'd8921 : data_rom <= {16'd24732, 16'd21495};
                15'd8922 : data_rom <= {16'd24734, 16'd21493};
                15'd8923 : data_rom <= {16'd24736, 16'd21491};
                15'd8924 : data_rom <= {16'd24738, 16'd21488};
                15'd8925 : data_rom <= {16'd24740, 16'd21486};
                15'd8926 : data_rom <= {16'd24742, 16'd21483};
                15'd8927 : data_rom <= {16'd24744, 16'd21481};
                15'd8928 : data_rom <= {16'd24746, 16'd21479};
                15'd8929 : data_rom <= {16'd24748, 16'd21476};
                15'd8930 : data_rom <= {16'd24750, 16'd21474};
                15'd8931 : data_rom <= {16'd24752, 16'd21472};
                15'd8932 : data_rom <= {16'd24754, 16'd21469};
                15'd8933 : data_rom <= {16'd24756, 16'd21467};
                15'd8934 : data_rom <= {16'd24758, 16'd21464};
                15'd8935 : data_rom <= {16'd24760, 16'd21462};
                15'd8936 : data_rom <= {16'd24762, 16'd21460};
                15'd8937 : data_rom <= {16'd24764, 16'd21457};
                15'd8938 : data_rom <= {16'd24767, 16'd21455};
                15'd8939 : data_rom <= {16'd24769, 16'd21453};
                15'd8940 : data_rom <= {16'd24771, 16'd21450};
                15'd8941 : data_rom <= {16'd24773, 16'd21448};
                15'd8942 : data_rom <= {16'd24775, 16'd21445};
                15'd8943 : data_rom <= {16'd24777, 16'd21443};
                15'd8944 : data_rom <= {16'd24779, 16'd21441};
                15'd8945 : data_rom <= {16'd24781, 16'd21438};
                15'd8946 : data_rom <= {16'd24783, 16'd21436};
                15'd8947 : data_rom <= {16'd24785, 16'd21434};
                15'd8948 : data_rom <= {16'd24787, 16'd21431};
                15'd8949 : data_rom <= {16'd24789, 16'd21429};
                15'd8950 : data_rom <= {16'd24791, 16'd21426};
                15'd8951 : data_rom <= {16'd24793, 16'd21424};
                15'd8952 : data_rom <= {16'd24795, 16'd21422};
                15'd8953 : data_rom <= {16'd24797, 16'd21419};
                15'd8954 : data_rom <= {16'd24799, 16'd21417};
                15'd8955 : data_rom <= {16'd24801, 16'd21415};
                15'd8956 : data_rom <= {16'd24803, 16'd21412};
                15'd8957 : data_rom <= {16'd24806, 16'd21410};
                15'd8958 : data_rom <= {16'd24808, 16'd21407};
                15'd8959 : data_rom <= {16'd24810, 16'd21405};
                15'd8960 : data_rom <= {16'd24812, 16'd21403};
                15'd8961 : data_rom <= {16'd24814, 16'd21400};
                15'd8962 : data_rom <= {16'd24816, 16'd21398};
                15'd8963 : data_rom <= {16'd24818, 16'd21396};
                15'd8964 : data_rom <= {16'd24820, 16'd21393};
                15'd8965 : data_rom <= {16'd24822, 16'd21391};
                15'd8966 : data_rom <= {16'd24824, 16'd21388};
                15'd8967 : data_rom <= {16'd24826, 16'd21386};
                15'd8968 : data_rom <= {16'd24828, 16'd21384};
                15'd8969 : data_rom <= {16'd24830, 16'd21381};
                15'd8970 : data_rom <= {16'd24832, 16'd21379};
                15'd8971 : data_rom <= {16'd24834, 16'd21377};
                15'd8972 : data_rom <= {16'd24836, 16'd21374};
                15'd8973 : data_rom <= {16'd24838, 16'd21372};
                15'd8974 : data_rom <= {16'd24840, 16'd21369};
                15'd8975 : data_rom <= {16'd24842, 16'd21367};
                15'd8976 : data_rom <= {16'd24845, 16'd21365};
                15'd8977 : data_rom <= {16'd24847, 16'd21362};
                15'd8978 : data_rom <= {16'd24849, 16'd21360};
                15'd8979 : data_rom <= {16'd24851, 16'd21357};
                15'd8980 : data_rom <= {16'd24853, 16'd21355};
                15'd8981 : data_rom <= {16'd24855, 16'd21353};
                15'd8982 : data_rom <= {16'd24857, 16'd21350};
                15'd8983 : data_rom <= {16'd24859, 16'd21348};
                15'd8984 : data_rom <= {16'd24861, 16'd21346};
                15'd8985 : data_rom <= {16'd24863, 16'd21343};
                15'd8986 : data_rom <= {16'd24865, 16'd21341};
                15'd8987 : data_rom <= {16'd24867, 16'd21338};
                15'd8988 : data_rom <= {16'd24869, 16'd21336};
                15'd8989 : data_rom <= {16'd24871, 16'd21334};
                15'd8990 : data_rom <= {16'd24873, 16'd21331};
                15'd8991 : data_rom <= {16'd24875, 16'd21329};
                15'd8992 : data_rom <= {16'd24877, 16'd21326};
                15'd8993 : data_rom <= {16'd24879, 16'd21324};
                15'd8994 : data_rom <= {16'd24881, 16'd21322};
                15'd8995 : data_rom <= {16'd24883, 16'd21319};
                15'd8996 : data_rom <= {16'd24885, 16'd21317};
                15'd8997 : data_rom <= {16'd24887, 16'd21315};
                15'd8998 : data_rom <= {16'd24890, 16'd21312};
                15'd8999 : data_rom <= {16'd24892, 16'd21310};
                15'd9000 : data_rom <= {16'd24894, 16'd21307};
                15'd9001 : data_rom <= {16'd24896, 16'd21305};
                15'd9002 : data_rom <= {16'd24898, 16'd21303};
                15'd9003 : data_rom <= {16'd24900, 16'd21300};
                15'd9004 : data_rom <= {16'd24902, 16'd21298};
                15'd9005 : data_rom <= {16'd24904, 16'd21295};
                15'd9006 : data_rom <= {16'd24906, 16'd21293};
                15'd9007 : data_rom <= {16'd24908, 16'd21291};
                15'd9008 : data_rom <= {16'd24910, 16'd21288};
                15'd9009 : data_rom <= {16'd24912, 16'd21286};
                15'd9010 : data_rom <= {16'd24914, 16'd21284};
                15'd9011 : data_rom <= {16'd24916, 16'd21281};
                15'd9012 : data_rom <= {16'd24918, 16'd21279};
                15'd9013 : data_rom <= {16'd24920, 16'd21276};
                15'd9014 : data_rom <= {16'd24922, 16'd21274};
                15'd9015 : data_rom <= {16'd24924, 16'd21272};
                15'd9016 : data_rom <= {16'd24926, 16'd21269};
                15'd9017 : data_rom <= {16'd24928, 16'd21267};
                15'd9018 : data_rom <= {16'd24930, 16'd21264};
                15'd9019 : data_rom <= {16'd24932, 16'd21262};
                15'd9020 : data_rom <= {16'd24934, 16'd21260};
                15'd9021 : data_rom <= {16'd24936, 16'd21257};
                15'd9022 : data_rom <= {16'd24938, 16'd21255};
                15'd9023 : data_rom <= {16'd24941, 16'd21252};
                15'd9024 : data_rom <= {16'd24943, 16'd21250};
                15'd9025 : data_rom <= {16'd24945, 16'd21248};
                15'd9026 : data_rom <= {16'd24947, 16'd21245};
                15'd9027 : data_rom <= {16'd24949, 16'd21243};
                15'd9028 : data_rom <= {16'd24951, 16'd21240};
                15'd9029 : data_rom <= {16'd24953, 16'd21238};
                15'd9030 : data_rom <= {16'd24955, 16'd21236};
                15'd9031 : data_rom <= {16'd24957, 16'd21233};
                15'd9032 : data_rom <= {16'd24959, 16'd21231};
                15'd9033 : data_rom <= {16'd24961, 16'd21229};
                15'd9034 : data_rom <= {16'd24963, 16'd21226};
                15'd9035 : data_rom <= {16'd24965, 16'd21224};
                15'd9036 : data_rom <= {16'd24967, 16'd21221};
                15'd9037 : data_rom <= {16'd24969, 16'd21219};
                15'd9038 : data_rom <= {16'd24971, 16'd21217};
                15'd9039 : data_rom <= {16'd24973, 16'd21214};
                15'd9040 : data_rom <= {16'd24975, 16'd21212};
                15'd9041 : data_rom <= {16'd24977, 16'd21209};
                15'd9042 : data_rom <= {16'd24979, 16'd21207};
                15'd9043 : data_rom <= {16'd24981, 16'd21205};
                15'd9044 : data_rom <= {16'd24983, 16'd21202};
                15'd9045 : data_rom <= {16'd24985, 16'd21200};
                15'd9046 : data_rom <= {16'd24987, 16'd21197};
                15'd9047 : data_rom <= {16'd24989, 16'd21195};
                15'd9048 : data_rom <= {16'd24991, 16'd21193};
                15'd9049 : data_rom <= {16'd24993, 16'd21190};
                15'd9050 : data_rom <= {16'd24995, 16'd21188};
                15'd9051 : data_rom <= {16'd24997, 16'd21185};
                15'd9052 : data_rom <= {16'd25000, 16'd21183};
                15'd9053 : data_rom <= {16'd25002, 16'd21181};
                15'd9054 : data_rom <= {16'd25004, 16'd21178};
                15'd9055 : data_rom <= {16'd25006, 16'd21176};
                15'd9056 : data_rom <= {16'd25008, 16'd21173};
                15'd9057 : data_rom <= {16'd25010, 16'd21171};
                15'd9058 : data_rom <= {16'd25012, 16'd21169};
                15'd9059 : data_rom <= {16'd25014, 16'd21166};
                15'd9060 : data_rom <= {16'd25016, 16'd21164};
                15'd9061 : data_rom <= {16'd25018, 16'd21161};
                15'd9062 : data_rom <= {16'd25020, 16'd21159};
                15'd9063 : data_rom <= {16'd25022, 16'd21157};
                15'd9064 : data_rom <= {16'd25024, 16'd21154};
                15'd9065 : data_rom <= {16'd25026, 16'd21152};
                15'd9066 : data_rom <= {16'd25028, 16'd21149};
                15'd9067 : data_rom <= {16'd25030, 16'd21147};
                15'd9068 : data_rom <= {16'd25032, 16'd21145};
                15'd9069 : data_rom <= {16'd25034, 16'd21142};
                15'd9070 : data_rom <= {16'd25036, 16'd21140};
                15'd9071 : data_rom <= {16'd25038, 16'd21137};
                15'd9072 : data_rom <= {16'd25040, 16'd21135};
                15'd9073 : data_rom <= {16'd25042, 16'd21133};
                15'd9074 : data_rom <= {16'd25044, 16'd21130};
                15'd9075 : data_rom <= {16'd25046, 16'd21128};
                15'd9076 : data_rom <= {16'd25048, 16'd21125};
                15'd9077 : data_rom <= {16'd25050, 16'd21123};
                15'd9078 : data_rom <= {16'd25052, 16'd21121};
                15'd9079 : data_rom <= {16'd25054, 16'd21118};
                15'd9080 : data_rom <= {16'd25056, 16'd21116};
                15'd9081 : data_rom <= {16'd25058, 16'd21113};
                15'd9082 : data_rom <= {16'd25060, 16'd21111};
                15'd9083 : data_rom <= {16'd25062, 16'd21109};
                15'd9084 : data_rom <= {16'd25064, 16'd21106};
                15'd9085 : data_rom <= {16'd25066, 16'd21104};
                15'd9086 : data_rom <= {16'd25068, 16'd21101};
                15'd9087 : data_rom <= {16'd25070, 16'd21099};
                15'd9088 : data_rom <= {16'd25072, 16'd21097};
                15'd9089 : data_rom <= {16'd25075, 16'd21094};
                15'd9090 : data_rom <= {16'd25077, 16'd21092};
                15'd9091 : data_rom <= {16'd25079, 16'd21089};
                15'd9092 : data_rom <= {16'd25081, 16'd21087};
                15'd9093 : data_rom <= {16'd25083, 16'd21085};
                15'd9094 : data_rom <= {16'd25085, 16'd21082};
                15'd9095 : data_rom <= {16'd25087, 16'd21080};
                15'd9096 : data_rom <= {16'd25089, 16'd21077};
                15'd9097 : data_rom <= {16'd25091, 16'd21075};
                15'd9098 : data_rom <= {16'd25093, 16'd21073};
                15'd9099 : data_rom <= {16'd25095, 16'd21070};
                15'd9100 : data_rom <= {16'd25097, 16'd21068};
                15'd9101 : data_rom <= {16'd25099, 16'd21065};
                15'd9102 : data_rom <= {16'd25101, 16'd21063};
                15'd9103 : data_rom <= {16'd25103, 16'd21061};
                15'd9104 : data_rom <= {16'd25105, 16'd21058};
                15'd9105 : data_rom <= {16'd25107, 16'd21056};
                15'd9106 : data_rom <= {16'd25109, 16'd21053};
                15'd9107 : data_rom <= {16'd25111, 16'd21051};
                15'd9108 : data_rom <= {16'd25113, 16'd21048};
                15'd9109 : data_rom <= {16'd25115, 16'd21046};
                15'd9110 : data_rom <= {16'd25117, 16'd21044};
                15'd9111 : data_rom <= {16'd25119, 16'd21041};
                15'd9112 : data_rom <= {16'd25121, 16'd21039};
                15'd9113 : data_rom <= {16'd25123, 16'd21036};
                15'd9114 : data_rom <= {16'd25125, 16'd21034};
                15'd9115 : data_rom <= {16'd25127, 16'd21032};
                15'd9116 : data_rom <= {16'd25129, 16'd21029};
                15'd9117 : data_rom <= {16'd25131, 16'd21027};
                15'd9118 : data_rom <= {16'd25133, 16'd21024};
                15'd9119 : data_rom <= {16'd25135, 16'd21022};
                15'd9120 : data_rom <= {16'd25137, 16'd21020};
                15'd9121 : data_rom <= {16'd25139, 16'd21017};
                15'd9122 : data_rom <= {16'd25141, 16'd21015};
                15'd9123 : data_rom <= {16'd25143, 16'd21012};
                15'd9124 : data_rom <= {16'd25145, 16'd21010};
                15'd9125 : data_rom <= {16'd25147, 16'd21008};
                15'd9126 : data_rom <= {16'd25149, 16'd21005};
                15'd9127 : data_rom <= {16'd25151, 16'd21003};
                15'd9128 : data_rom <= {16'd25153, 16'd21000};
                15'd9129 : data_rom <= {16'd25155, 16'd20998};
                15'd9130 : data_rom <= {16'd25157, 16'd20995};
                15'd9131 : data_rom <= {16'd25159, 16'd20993};
                15'd9132 : data_rom <= {16'd25161, 16'd20991};
                15'd9133 : data_rom <= {16'd25163, 16'd20988};
                15'd9134 : data_rom <= {16'd25165, 16'd20986};
                15'd9135 : data_rom <= {16'd25167, 16'd20983};
                15'd9136 : data_rom <= {16'd25169, 16'd20981};
                15'd9137 : data_rom <= {16'd25171, 16'd20979};
                15'd9138 : data_rom <= {16'd25173, 16'd20976};
                15'd9139 : data_rom <= {16'd25175, 16'd20974};
                15'd9140 : data_rom <= {16'd25177, 16'd20971};
                15'd9141 : data_rom <= {16'd25179, 16'd20969};
                15'd9142 : data_rom <= {16'd25181, 16'd20967};
                15'd9143 : data_rom <= {16'd25183, 16'd20964};
                15'd9144 : data_rom <= {16'd25185, 16'd20962};
                15'd9145 : data_rom <= {16'd25187, 16'd20959};
                15'd9146 : data_rom <= {16'd25189, 16'd20957};
                15'd9147 : data_rom <= {16'd25191, 16'd20954};
                15'd9148 : data_rom <= {16'd25193, 16'd20952};
                15'd9149 : data_rom <= {16'd25195, 16'd20950};
                15'd9150 : data_rom <= {16'd25197, 16'd20947};
                15'd9151 : data_rom <= {16'd25199, 16'd20945};
                15'd9152 : data_rom <= {16'd25201, 16'd20942};
                15'd9153 : data_rom <= {16'd25203, 16'd20940};
                15'd9154 : data_rom <= {16'd25205, 16'd20938};
                15'd9155 : data_rom <= {16'd25207, 16'd20935};
                15'd9156 : data_rom <= {16'd25209, 16'd20933};
                15'd9157 : data_rom <= {16'd25211, 16'd20930};
                15'd9158 : data_rom <= {16'd25214, 16'd20928};
                15'd9159 : data_rom <= {16'd25216, 16'd20925};
                15'd9160 : data_rom <= {16'd25218, 16'd20923};
                15'd9161 : data_rom <= {16'd25220, 16'd20921};
                15'd9162 : data_rom <= {16'd25222, 16'd20918};
                15'd9163 : data_rom <= {16'd25224, 16'd20916};
                15'd9164 : data_rom <= {16'd25226, 16'd20913};
                15'd9165 : data_rom <= {16'd25228, 16'd20911};
                15'd9166 : data_rom <= {16'd25230, 16'd20909};
                15'd9167 : data_rom <= {16'd25232, 16'd20906};
                15'd9168 : data_rom <= {16'd25234, 16'd20904};
                15'd9169 : data_rom <= {16'd25236, 16'd20901};
                15'd9170 : data_rom <= {16'd25238, 16'd20899};
                15'd9171 : data_rom <= {16'd25240, 16'd20896};
                15'd9172 : data_rom <= {16'd25242, 16'd20894};
                15'd9173 : data_rom <= {16'd25244, 16'd20892};
                15'd9174 : data_rom <= {16'd25246, 16'd20889};
                15'd9175 : data_rom <= {16'd25248, 16'd20887};
                15'd9176 : data_rom <= {16'd25250, 16'd20884};
                15'd9177 : data_rom <= {16'd25252, 16'd20882};
                15'd9178 : data_rom <= {16'd25254, 16'd20879};
                15'd9179 : data_rom <= {16'd25256, 16'd20877};
                15'd9180 : data_rom <= {16'd25258, 16'd20875};
                15'd9181 : data_rom <= {16'd25260, 16'd20872};
                15'd9182 : data_rom <= {16'd25262, 16'd20870};
                15'd9183 : data_rom <= {16'd25264, 16'd20867};
                15'd9184 : data_rom <= {16'd25266, 16'd20865};
                15'd9185 : data_rom <= {16'd25268, 16'd20863};
                15'd9186 : data_rom <= {16'd25270, 16'd20860};
                15'd9187 : data_rom <= {16'd25272, 16'd20858};
                15'd9188 : data_rom <= {16'd25274, 16'd20855};
                15'd9189 : data_rom <= {16'd25276, 16'd20853};
                15'd9190 : data_rom <= {16'd25278, 16'd20850};
                15'd9191 : data_rom <= {16'd25280, 16'd20848};
                15'd9192 : data_rom <= {16'd25282, 16'd20846};
                15'd9193 : data_rom <= {16'd25284, 16'd20843};
                15'd9194 : data_rom <= {16'd25286, 16'd20841};
                15'd9195 : data_rom <= {16'd25288, 16'd20838};
                15'd9196 : data_rom <= {16'd25290, 16'd20836};
                15'd9197 : data_rom <= {16'd25292, 16'd20833};
                15'd9198 : data_rom <= {16'd25294, 16'd20831};
                15'd9199 : data_rom <= {16'd25296, 16'd20829};
                15'd9200 : data_rom <= {16'd25298, 16'd20826};
                15'd9201 : data_rom <= {16'd25300, 16'd20824};
                15'd9202 : data_rom <= {16'd25302, 16'd20821};
                15'd9203 : data_rom <= {16'd25304, 16'd20819};
                15'd9204 : data_rom <= {16'd25306, 16'd20816};
                15'd9205 : data_rom <= {16'd25308, 16'd20814};
                15'd9206 : data_rom <= {16'd25310, 16'd20812};
                15'd9207 : data_rom <= {16'd25312, 16'd20809};
                15'd9208 : data_rom <= {16'd25314, 16'd20807};
                15'd9209 : data_rom <= {16'd25316, 16'd20804};
                15'd9210 : data_rom <= {16'd25318, 16'd20802};
                15'd9211 : data_rom <= {16'd25320, 16'd20799};
                15'd9212 : data_rom <= {16'd25322, 16'd20797};
                15'd9213 : data_rom <= {16'd25324, 16'd20795};
                15'd9214 : data_rom <= {16'd25326, 16'd20792};
                15'd9215 : data_rom <= {16'd25327, 16'd20790};
                15'd9216 : data_rom <= {16'd25329, 16'd20787};
                15'd9217 : data_rom <= {16'd25331, 16'd20785};
                15'd9218 : data_rom <= {16'd25333, 16'd20782};
                15'd9219 : data_rom <= {16'd25335, 16'd20780};
                15'd9220 : data_rom <= {16'd25337, 16'd20778};
                15'd9221 : data_rom <= {16'd25339, 16'd20775};
                15'd9222 : data_rom <= {16'd25341, 16'd20773};
                15'd9223 : data_rom <= {16'd25343, 16'd20770};
                15'd9224 : data_rom <= {16'd25345, 16'd20768};
                15'd9225 : data_rom <= {16'd25347, 16'd20765};
                15'd9226 : data_rom <= {16'd25349, 16'd20763};
                15'd9227 : data_rom <= {16'd25351, 16'd20761};
                15'd9228 : data_rom <= {16'd25353, 16'd20758};
                15'd9229 : data_rom <= {16'd25355, 16'd20756};
                15'd9230 : data_rom <= {16'd25357, 16'd20753};
                15'd9231 : data_rom <= {16'd25359, 16'd20751};
                15'd9232 : data_rom <= {16'd25361, 16'd20748};
                15'd9233 : data_rom <= {16'd25363, 16'd20746};
                15'd9234 : data_rom <= {16'd25365, 16'd20744};
                15'd9235 : data_rom <= {16'd25367, 16'd20741};
                15'd9236 : data_rom <= {16'd25369, 16'd20739};
                15'd9237 : data_rom <= {16'd25371, 16'd20736};
                15'd9238 : data_rom <= {16'd25373, 16'd20734};
                15'd9239 : data_rom <= {16'd25375, 16'd20731};
                15'd9240 : data_rom <= {16'd25377, 16'd20729};
                15'd9241 : data_rom <= {16'd25379, 16'd20727};
                15'd9242 : data_rom <= {16'd25381, 16'd20724};
                15'd9243 : data_rom <= {16'd25383, 16'd20722};
                15'd9244 : data_rom <= {16'd25385, 16'd20719};
                15'd9245 : data_rom <= {16'd25387, 16'd20717};
                15'd9246 : data_rom <= {16'd25389, 16'd20714};
                15'd9247 : data_rom <= {16'd25391, 16'd20712};
                15'd9248 : data_rom <= {16'd25393, 16'd20710};
                15'd9249 : data_rom <= {16'd25395, 16'd20707};
                15'd9250 : data_rom <= {16'd25397, 16'd20705};
                15'd9251 : data_rom <= {16'd25399, 16'd20702};
                15'd9252 : data_rom <= {16'd25401, 16'd20700};
                15'd9253 : data_rom <= {16'd25403, 16'd20697};
                15'd9254 : data_rom <= {16'd25405, 16'd20695};
                15'd9255 : data_rom <= {16'd25407, 16'd20692};
                15'd9256 : data_rom <= {16'd25409, 16'd20690};
                15'd9257 : data_rom <= {16'd25411, 16'd20688};
                15'd9258 : data_rom <= {16'd25413, 16'd20685};
                15'd9259 : data_rom <= {16'd25415, 16'd20683};
                15'd9260 : data_rom <= {16'd25417, 16'd20680};
                15'd9261 : data_rom <= {16'd25419, 16'd20678};
                15'd9262 : data_rom <= {16'd25421, 16'd20675};
                15'd9263 : data_rom <= {16'd25423, 16'd20673};
                15'd9264 : data_rom <= {16'd25425, 16'd20671};
                15'd9265 : data_rom <= {16'd25427, 16'd20668};
                15'd9266 : data_rom <= {16'd25429, 16'd20666};
                15'd9267 : data_rom <= {16'd25431, 16'd20663};
                15'd9268 : data_rom <= {16'd25433, 16'd20661};
                15'd9269 : data_rom <= {16'd25435, 16'd20658};
                15'd9270 : data_rom <= {16'd25437, 16'd20656};
                15'd9271 : data_rom <= {16'd25439, 16'd20653};
                15'd9272 : data_rom <= {16'd25441, 16'd20651};
                15'd9273 : data_rom <= {16'd25443, 16'd20649};
                15'd9274 : data_rom <= {16'd25445, 16'd20646};
                15'd9275 : data_rom <= {16'd25447, 16'd20644};
                15'd9276 : data_rom <= {16'd25449, 16'd20641};
                15'd9277 : data_rom <= {16'd25451, 16'd20639};
                15'd9278 : data_rom <= {16'd25453, 16'd20636};
                15'd9279 : data_rom <= {16'd25455, 16'd20634};
                15'd9280 : data_rom <= {16'd25457, 16'd20632};
                15'd9281 : data_rom <= {16'd25459, 16'd20629};
                15'd9282 : data_rom <= {16'd25461, 16'd20627};
                15'd9283 : data_rom <= {16'd25462, 16'd20624};
                15'd9284 : data_rom <= {16'd25464, 16'd20622};
                15'd9285 : data_rom <= {16'd25466, 16'd20619};
                15'd9286 : data_rom <= {16'd25468, 16'd20617};
                15'd9287 : data_rom <= {16'd25470, 16'd20614};
                15'd9288 : data_rom <= {16'd25472, 16'd20612};
                15'd9289 : data_rom <= {16'd25474, 16'd20610};
                15'd9290 : data_rom <= {16'd25476, 16'd20607};
                15'd9291 : data_rom <= {16'd25478, 16'd20605};
                15'd9292 : data_rom <= {16'd25480, 16'd20602};
                15'd9293 : data_rom <= {16'd25482, 16'd20600};
                15'd9294 : data_rom <= {16'd25484, 16'd20597};
                15'd9295 : data_rom <= {16'd25486, 16'd20595};
                15'd9296 : data_rom <= {16'd25488, 16'd20592};
                15'd9297 : data_rom <= {16'd25490, 16'd20590};
                15'd9298 : data_rom <= {16'd25492, 16'd20588};
                15'd9299 : data_rom <= {16'd25494, 16'd20585};
                15'd9300 : data_rom <= {16'd25496, 16'd20583};
                15'd9301 : data_rom <= {16'd25498, 16'd20580};
                15'd9302 : data_rom <= {16'd25500, 16'd20578};
                15'd9303 : data_rom <= {16'd25502, 16'd20575};
                15'd9304 : data_rom <= {16'd25504, 16'd20573};
                15'd9305 : data_rom <= {16'd25506, 16'd20570};
                15'd9306 : data_rom <= {16'd25508, 16'd20568};
                15'd9307 : data_rom <= {16'd25510, 16'd20566};
                15'd9308 : data_rom <= {16'd25512, 16'd20563};
                15'd9309 : data_rom <= {16'd25514, 16'd20561};
                15'd9310 : data_rom <= {16'd25516, 16'd20558};
                15'd9311 : data_rom <= {16'd25518, 16'd20556};
                15'd9312 : data_rom <= {16'd25520, 16'd20553};
                15'd9313 : data_rom <= {16'd25522, 16'd20551};
                15'd9314 : data_rom <= {16'd25524, 16'd20548};
                15'd9315 : data_rom <= {16'd25526, 16'd20546};
                15'd9316 : data_rom <= {16'd25528, 16'd20544};
                15'd9317 : data_rom <= {16'd25530, 16'd20541};
                15'd9318 : data_rom <= {16'd25532, 16'd20539};
                15'd9319 : data_rom <= {16'd25534, 16'd20536};
                15'd9320 : data_rom <= {16'd25535, 16'd20534};
                15'd9321 : data_rom <= {16'd25537, 16'd20531};
                15'd9322 : data_rom <= {16'd25539, 16'd20529};
                15'd9323 : data_rom <= {16'd25541, 16'd20526};
                15'd9324 : data_rom <= {16'd25543, 16'd20524};
                15'd9325 : data_rom <= {16'd25545, 16'd20521};
                15'd9326 : data_rom <= {16'd25547, 16'd20519};
                15'd9327 : data_rom <= {16'd25549, 16'd20517};
                15'd9328 : data_rom <= {16'd25551, 16'd20514};
                15'd9329 : data_rom <= {16'd25553, 16'd20512};
                15'd9330 : data_rom <= {16'd25555, 16'd20509};
                15'd9331 : data_rom <= {16'd25557, 16'd20507};
                15'd9332 : data_rom <= {16'd25559, 16'd20504};
                15'd9333 : data_rom <= {16'd25561, 16'd20502};
                15'd9334 : data_rom <= {16'd25563, 16'd20499};
                15'd9335 : data_rom <= {16'd25565, 16'd20497};
                15'd9336 : data_rom <= {16'd25567, 16'd20495};
                15'd9337 : data_rom <= {16'd25569, 16'd20492};
                15'd9338 : data_rom <= {16'd25571, 16'd20490};
                15'd9339 : data_rom <= {16'd25573, 16'd20487};
                15'd9340 : data_rom <= {16'd25575, 16'd20485};
                15'd9341 : data_rom <= {16'd25577, 16'd20482};
                15'd9342 : data_rom <= {16'd25579, 16'd20480};
                15'd9343 : data_rom <= {16'd25581, 16'd20477};
                15'd9344 : data_rom <= {16'd25583, 16'd20475};
                15'd9345 : data_rom <= {16'd25585, 16'd20472};
                15'd9346 : data_rom <= {16'd25587, 16'd20470};
                15'd9347 : data_rom <= {16'd25589, 16'd20468};
                15'd9348 : data_rom <= {16'd25591, 16'd20465};
                15'd9349 : data_rom <= {16'd25592, 16'd20463};
                15'd9350 : data_rom <= {16'd25594, 16'd20460};
                15'd9351 : data_rom <= {16'd25596, 16'd20458};
                15'd9352 : data_rom <= {16'd25598, 16'd20455};
                15'd9353 : data_rom <= {16'd25600, 16'd20453};
                15'd9354 : data_rom <= {16'd25602, 16'd20450};
                15'd9355 : data_rom <= {16'd25604, 16'd20448};
                15'd9356 : data_rom <= {16'd25606, 16'd20445};
                15'd9357 : data_rom <= {16'd25608, 16'd20443};
                15'd9358 : data_rom <= {16'd25610, 16'd20441};
                15'd9359 : data_rom <= {16'd25612, 16'd20438};
                15'd9360 : data_rom <= {16'd25614, 16'd20436};
                15'd9361 : data_rom <= {16'd25616, 16'd20433};
                15'd9362 : data_rom <= {16'd25618, 16'd20431};
                15'd9363 : data_rom <= {16'd25620, 16'd20428};
                15'd9364 : data_rom <= {16'd25622, 16'd20426};
                15'd9365 : data_rom <= {16'd25624, 16'd20423};
                15'd9366 : data_rom <= {16'd25626, 16'd20421};
                15'd9367 : data_rom <= {16'd25628, 16'd20418};
                15'd9368 : data_rom <= {16'd25630, 16'd20416};
                15'd9369 : data_rom <= {16'd25632, 16'd20414};
                15'd9370 : data_rom <= {16'd25634, 16'd20411};
                15'd9371 : data_rom <= {16'd25636, 16'd20409};
                15'd9372 : data_rom <= {16'd25638, 16'd20406};
                15'd9373 : data_rom <= {16'd25640, 16'd20404};
                15'd9374 : data_rom <= {16'd25641, 16'd20401};
                15'd9375 : data_rom <= {16'd25643, 16'd20399};
                15'd9376 : data_rom <= {16'd25645, 16'd20396};
                15'd9377 : data_rom <= {16'd25647, 16'd20394};
                15'd9378 : data_rom <= {16'd25649, 16'd20391};
                15'd9379 : data_rom <= {16'd25651, 16'd20389};
                15'd9380 : data_rom <= {16'd25653, 16'd20386};
                15'd9381 : data_rom <= {16'd25655, 16'd20384};
                15'd9382 : data_rom <= {16'd25657, 16'd20382};
                15'd9383 : data_rom <= {16'd25659, 16'd20379};
                15'd9384 : data_rom <= {16'd25661, 16'd20377};
                15'd9385 : data_rom <= {16'd25663, 16'd20374};
                15'd9386 : data_rom <= {16'd25665, 16'd20372};
                15'd9387 : data_rom <= {16'd25667, 16'd20369};
                15'd9388 : data_rom <= {16'd25669, 16'd20367};
                15'd9389 : data_rom <= {16'd25671, 16'd20364};
                15'd9390 : data_rom <= {16'd25673, 16'd20362};
                15'd9391 : data_rom <= {16'd25675, 16'd20359};
                15'd9392 : data_rom <= {16'd25677, 16'd20357};
                15'd9393 : data_rom <= {16'd25679, 16'd20355};
                15'd9394 : data_rom <= {16'd25681, 16'd20352};
                15'd9395 : data_rom <= {16'd25682, 16'd20350};
                15'd9396 : data_rom <= {16'd25684, 16'd20347};
                15'd9397 : data_rom <= {16'd25686, 16'd20345};
                15'd9398 : data_rom <= {16'd25688, 16'd20342};
                15'd9399 : data_rom <= {16'd25690, 16'd20340};
                15'd9400 : data_rom <= {16'd25692, 16'd20337};
                15'd9401 : data_rom <= {16'd25694, 16'd20335};
                15'd9402 : data_rom <= {16'd25696, 16'd20332};
                15'd9403 : data_rom <= {16'd25698, 16'd20330};
                15'd9404 : data_rom <= {16'd25700, 16'd20327};
                15'd9405 : data_rom <= {16'd25702, 16'd20325};
                15'd9406 : data_rom <= {16'd25704, 16'd20322};
                15'd9407 : data_rom <= {16'd25706, 16'd20320};
                15'd9408 : data_rom <= {16'd25708, 16'd20318};
                15'd9409 : data_rom <= {16'd25710, 16'd20315};
                15'd9410 : data_rom <= {16'd25712, 16'd20313};
                15'd9411 : data_rom <= {16'd25714, 16'd20310};
                15'd9412 : data_rom <= {16'd25716, 16'd20308};
                15'd9413 : data_rom <= {16'd25718, 16'd20305};
                15'd9414 : data_rom <= {16'd25720, 16'd20303};
                15'd9415 : data_rom <= {16'd25721, 16'd20300};
                15'd9416 : data_rom <= {16'd25723, 16'd20298};
                15'd9417 : data_rom <= {16'd25725, 16'd20295};
                15'd9418 : data_rom <= {16'd25727, 16'd20293};
                15'd9419 : data_rom <= {16'd25729, 16'd20290};
                15'd9420 : data_rom <= {16'd25731, 16'd20288};
                15'd9421 : data_rom <= {16'd25733, 16'd20285};
                15'd9422 : data_rom <= {16'd25735, 16'd20283};
                15'd9423 : data_rom <= {16'd25737, 16'd20281};
                15'd9424 : data_rom <= {16'd25739, 16'd20278};
                15'd9425 : data_rom <= {16'd25741, 16'd20276};
                15'd9426 : data_rom <= {16'd25743, 16'd20273};
                15'd9427 : data_rom <= {16'd25745, 16'd20271};
                15'd9428 : data_rom <= {16'd25747, 16'd20268};
                15'd9429 : data_rom <= {16'd25749, 16'd20266};
                15'd9430 : data_rom <= {16'd25751, 16'd20263};
                15'd9431 : data_rom <= {16'd25753, 16'd20261};
                15'd9432 : data_rom <= {16'd25755, 16'd20258};
                15'd9433 : data_rom <= {16'd25756, 16'd20256};
                15'd9434 : data_rom <= {16'd25758, 16'd20253};
                15'd9435 : data_rom <= {16'd25760, 16'd20251};
                15'd9436 : data_rom <= {16'd25762, 16'd20248};
                15'd9437 : data_rom <= {16'd25764, 16'd20246};
                15'd9438 : data_rom <= {16'd25766, 16'd20244};
                15'd9439 : data_rom <= {16'd25768, 16'd20241};
                15'd9440 : data_rom <= {16'd25770, 16'd20239};
                15'd9441 : data_rom <= {16'd25772, 16'd20236};
                15'd9442 : data_rom <= {16'd25774, 16'd20234};
                15'd9443 : data_rom <= {16'd25776, 16'd20231};
                15'd9444 : data_rom <= {16'd25778, 16'd20229};
                15'd9445 : data_rom <= {16'd25780, 16'd20226};
                15'd9446 : data_rom <= {16'd25782, 16'd20224};
                15'd9447 : data_rom <= {16'd25784, 16'd20221};
                15'd9448 : data_rom <= {16'd25786, 16'd20219};
                15'd9449 : data_rom <= {16'd25788, 16'd20216};
                15'd9450 : data_rom <= {16'd25789, 16'd20214};
                15'd9451 : data_rom <= {16'd25791, 16'd20211};
                15'd9452 : data_rom <= {16'd25793, 16'd20209};
                15'd9453 : data_rom <= {16'd25795, 16'd20206};
                15'd9454 : data_rom <= {16'd25797, 16'd20204};
                15'd9455 : data_rom <= {16'd25799, 16'd20202};
                15'd9456 : data_rom <= {16'd25801, 16'd20199};
                15'd9457 : data_rom <= {16'd25803, 16'd20197};
                15'd9458 : data_rom <= {16'd25805, 16'd20194};
                15'd9459 : data_rom <= {16'd25807, 16'd20192};
                15'd9460 : data_rom <= {16'd25809, 16'd20189};
                15'd9461 : data_rom <= {16'd25811, 16'd20187};
                15'd9462 : data_rom <= {16'd25813, 16'd20184};
                15'd9463 : data_rom <= {16'd25815, 16'd20182};
                15'd9464 : data_rom <= {16'd25817, 16'd20179};
                15'd9465 : data_rom <= {16'd25818, 16'd20177};
                15'd9466 : data_rom <= {16'd25820, 16'd20174};
                15'd9467 : data_rom <= {16'd25822, 16'd20172};
                15'd9468 : data_rom <= {16'd25824, 16'd20169};
                15'd9469 : data_rom <= {16'd25826, 16'd20167};
                15'd9470 : data_rom <= {16'd25828, 16'd20164};
                15'd9471 : data_rom <= {16'd25830, 16'd20162};
                15'd9472 : data_rom <= {16'd25832, 16'd20159};
                15'd9473 : data_rom <= {16'd25834, 16'd20157};
                15'd9474 : data_rom <= {16'd25836, 16'd20154};
                15'd9475 : data_rom <= {16'd25838, 16'd20152};
                15'd9476 : data_rom <= {16'd25840, 16'd20150};
                15'd9477 : data_rom <= {16'd25842, 16'd20147};
                15'd9478 : data_rom <= {16'd25844, 16'd20145};
                15'd9479 : data_rom <= {16'd25846, 16'd20142};
                15'd9480 : data_rom <= {16'd25847, 16'd20140};
                15'd9481 : data_rom <= {16'd25849, 16'd20137};
                15'd9482 : data_rom <= {16'd25851, 16'd20135};
                15'd9483 : data_rom <= {16'd25853, 16'd20132};
                15'd9484 : data_rom <= {16'd25855, 16'd20130};
                15'd9485 : data_rom <= {16'd25857, 16'd20127};
                15'd9486 : data_rom <= {16'd25859, 16'd20125};
                15'd9487 : data_rom <= {16'd25861, 16'd20122};
                15'd9488 : data_rom <= {16'd25863, 16'd20120};
                15'd9489 : data_rom <= {16'd25865, 16'd20117};
                15'd9490 : data_rom <= {16'd25867, 16'd20115};
                15'd9491 : data_rom <= {16'd25869, 16'd20112};
                15'd9492 : data_rom <= {16'd25871, 16'd20110};
                15'd9493 : data_rom <= {16'd25873, 16'd20107};
                15'd9494 : data_rom <= {16'd25874, 16'd20105};
                15'd9495 : data_rom <= {16'd25876, 16'd20102};
                15'd9496 : data_rom <= {16'd25878, 16'd20100};
                15'd9497 : data_rom <= {16'd25880, 16'd20097};
                15'd9498 : data_rom <= {16'd25882, 16'd20095};
                15'd9499 : data_rom <= {16'd25884, 16'd20092};
                15'd9500 : data_rom <= {16'd25886, 16'd20090};
                15'd9501 : data_rom <= {16'd25888, 16'd20088};
                15'd9502 : data_rom <= {16'd25890, 16'd20085};
                15'd9503 : data_rom <= {16'd25892, 16'd20083};
                15'd9504 : data_rom <= {16'd25894, 16'd20080};
                15'd9505 : data_rom <= {16'd25896, 16'd20078};
                15'd9506 : data_rom <= {16'd25898, 16'd20075};
                15'd9507 : data_rom <= {16'd25900, 16'd20073};
                15'd9508 : data_rom <= {16'd25901, 16'd20070};
                15'd9509 : data_rom <= {16'd25903, 16'd20068};
                15'd9510 : data_rom <= {16'd25905, 16'd20065};
                15'd9511 : data_rom <= {16'd25907, 16'd20063};
                15'd9512 : data_rom <= {16'd25909, 16'd20060};
                15'd9513 : data_rom <= {16'd25911, 16'd20058};
                15'd9514 : data_rom <= {16'd25913, 16'd20055};
                15'd9515 : data_rom <= {16'd25915, 16'd20053};
                15'd9516 : data_rom <= {16'd25917, 16'd20050};
                15'd9517 : data_rom <= {16'd25919, 16'd20048};
                15'd9518 : data_rom <= {16'd25921, 16'd20045};
                15'd9519 : data_rom <= {16'd25923, 16'd20043};
                15'd9520 : data_rom <= {16'd25925, 16'd20040};
                15'd9521 : data_rom <= {16'd25926, 16'd20038};
                15'd9522 : data_rom <= {16'd25928, 16'd20035};
                15'd9523 : data_rom <= {16'd25930, 16'd20033};
                15'd9524 : data_rom <= {16'd25932, 16'd20030};
                15'd9525 : data_rom <= {16'd25934, 16'd20028};
                15'd9526 : data_rom <= {16'd25936, 16'd20025};
                15'd9527 : data_rom <= {16'd25938, 16'd20023};
                15'd9528 : data_rom <= {16'd25940, 16'd20020};
                15'd9529 : data_rom <= {16'd25942, 16'd20018};
                15'd9530 : data_rom <= {16'd25944, 16'd20015};
                15'd9531 : data_rom <= {16'd25946, 16'd20013};
                15'd9532 : data_rom <= {16'd25948, 16'd20010};
                15'd9533 : data_rom <= {16'd25949, 16'd20008};
                15'd9534 : data_rom <= {16'd25951, 16'd20006};
                15'd9535 : data_rom <= {16'd25953, 16'd20003};
                15'd9536 : data_rom <= {16'd25955, 16'd20001};
                15'd9537 : data_rom <= {16'd25957, 16'd19998};
                15'd9538 : data_rom <= {16'd25959, 16'd19996};
                15'd9539 : data_rom <= {16'd25961, 16'd19993};
                15'd9540 : data_rom <= {16'd25963, 16'd19991};
                15'd9541 : data_rom <= {16'd25965, 16'd19988};
                15'd9542 : data_rom <= {16'd25967, 16'd19986};
                15'd9543 : data_rom <= {16'd25969, 16'd19983};
                15'd9544 : data_rom <= {16'd25971, 16'd19981};
                15'd9545 : data_rom <= {16'd25972, 16'd19978};
                15'd9546 : data_rom <= {16'd25974, 16'd19976};
                15'd9547 : data_rom <= {16'd25976, 16'd19973};
                15'd9548 : data_rom <= {16'd25978, 16'd19971};
                15'd9549 : data_rom <= {16'd25980, 16'd19968};
                15'd9550 : data_rom <= {16'd25982, 16'd19966};
                15'd9551 : data_rom <= {16'd25984, 16'd19963};
                15'd9552 : data_rom <= {16'd25986, 16'd19961};
                15'd9553 : data_rom <= {16'd25988, 16'd19958};
                15'd9554 : data_rom <= {16'd25990, 16'd19956};
                15'd9555 : data_rom <= {16'd25992, 16'd19953};
                15'd9556 : data_rom <= {16'd25994, 16'd19951};
                15'd9557 : data_rom <= {16'd25995, 16'd19948};
                15'd9558 : data_rom <= {16'd25997, 16'd19946};
                15'd9559 : data_rom <= {16'd25999, 16'd19943};
                15'd9560 : data_rom <= {16'd26001, 16'd19941};
                15'd9561 : data_rom <= {16'd26003, 16'd19938};
                15'd9562 : data_rom <= {16'd26005, 16'd19936};
                15'd9563 : data_rom <= {16'd26007, 16'd19933};
                15'd9564 : data_rom <= {16'd26009, 16'd19931};
                15'd9565 : data_rom <= {16'd26011, 16'd19928};
                15'd9566 : data_rom <= {16'd26013, 16'd19926};
                15'd9567 : data_rom <= {16'd26015, 16'd19923};
                15'd9568 : data_rom <= {16'd26016, 16'd19921};
                15'd9569 : data_rom <= {16'd26018, 16'd19918};
                15'd9570 : data_rom <= {16'd26020, 16'd19916};
                15'd9571 : data_rom <= {16'd26022, 16'd19913};
                15'd9572 : data_rom <= {16'd26024, 16'd19911};
                15'd9573 : data_rom <= {16'd26026, 16'd19908};
                15'd9574 : data_rom <= {16'd26028, 16'd19906};
                15'd9575 : data_rom <= {16'd26030, 16'd19903};
                15'd9576 : data_rom <= {16'd26032, 16'd19901};
                15'd9577 : data_rom <= {16'd26034, 16'd19898};
                15'd9578 : data_rom <= {16'd26036, 16'd19896};
                15'd9579 : data_rom <= {16'd26037, 16'd19893};
                15'd9580 : data_rom <= {16'd26039, 16'd19891};
                15'd9581 : data_rom <= {16'd26041, 16'd19888};
                15'd9582 : data_rom <= {16'd26043, 16'd19886};
                15'd9583 : data_rom <= {16'd26045, 16'd19883};
                15'd9584 : data_rom <= {16'd26047, 16'd19881};
                15'd9585 : data_rom <= {16'd26049, 16'd19878};
                15'd9586 : data_rom <= {16'd26051, 16'd19876};
                15'd9587 : data_rom <= {16'd26053, 16'd19873};
                15'd9588 : data_rom <= {16'd26055, 16'd19871};
                15'd9589 : data_rom <= {16'd26057, 16'd19868};
                15'd9590 : data_rom <= {16'd26058, 16'd19866};
                15'd9591 : data_rom <= {16'd26060, 16'd19863};
                15'd9592 : data_rom <= {16'd26062, 16'd19861};
                15'd9593 : data_rom <= {16'd26064, 16'd19858};
                15'd9594 : data_rom <= {16'd26066, 16'd19856};
                15'd9595 : data_rom <= {16'd26068, 16'd19853};
                15'd9596 : data_rom <= {16'd26070, 16'd19851};
                15'd9597 : data_rom <= {16'd26072, 16'd19848};
                15'd9598 : data_rom <= {16'd26074, 16'd19846};
                15'd9599 : data_rom <= {16'd26076, 16'd19843};
                15'd9600 : data_rom <= {16'd26077, 16'd19841};
                15'd9601 : data_rom <= {16'd26079, 16'd19838};
                15'd9602 : data_rom <= {16'd26081, 16'd19836};
                15'd9603 : data_rom <= {16'd26083, 16'd19833};
                15'd9604 : data_rom <= {16'd26085, 16'd19831};
                15'd9605 : data_rom <= {16'd26087, 16'd19828};
                15'd9606 : data_rom <= {16'd26089, 16'd19826};
                15'd9607 : data_rom <= {16'd26091, 16'd19823};
                15'd9608 : data_rom <= {16'd26093, 16'd19821};
                15'd9609 : data_rom <= {16'd26095, 16'd19818};
                15'd9610 : data_rom <= {16'd26096, 16'd19816};
                15'd9611 : data_rom <= {16'd26098, 16'd19813};
                15'd9612 : data_rom <= {16'd26100, 16'd19811};
                15'd9613 : data_rom <= {16'd26102, 16'd19808};
                15'd9614 : data_rom <= {16'd26104, 16'd19806};
                15'd9615 : data_rom <= {16'd26106, 16'd19803};
                15'd9616 : data_rom <= {16'd26108, 16'd19801};
                15'd9617 : data_rom <= {16'd26110, 16'd19798};
                15'd9618 : data_rom <= {16'd26112, 16'd19796};
                15'd9619 : data_rom <= {16'd26114, 16'd19793};
                15'd9620 : data_rom <= {16'd26115, 16'd19791};
                15'd9621 : data_rom <= {16'd26117, 16'd19788};
                15'd9622 : data_rom <= {16'd26119, 16'd19786};
                15'd9623 : data_rom <= {16'd26121, 16'd19783};
                15'd9624 : data_rom <= {16'd26123, 16'd19781};
                15'd9625 : data_rom <= {16'd26125, 16'd19778};
                15'd9626 : data_rom <= {16'd26127, 16'd19776};
                15'd9627 : data_rom <= {16'd26129, 16'd19773};
                15'd9628 : data_rom <= {16'd26131, 16'd19771};
                15'd9629 : data_rom <= {16'd26133, 16'd19768};
                15'd9630 : data_rom <= {16'd26134, 16'd19766};
                15'd9631 : data_rom <= {16'd26136, 16'd19763};
                15'd9632 : data_rom <= {16'd26138, 16'd19761};
                15'd9633 : data_rom <= {16'd26140, 16'd19758};
                15'd9634 : data_rom <= {16'd26142, 16'd19756};
                15'd9635 : data_rom <= {16'd26144, 16'd19753};
                15'd9636 : data_rom <= {16'd26146, 16'd19751};
                15'd9637 : data_rom <= {16'd26148, 16'd19748};
                15'd9638 : data_rom <= {16'd26150, 16'd19746};
                15'd9639 : data_rom <= {16'd26151, 16'd19743};
                15'd9640 : data_rom <= {16'd26153, 16'd19741};
                15'd9641 : data_rom <= {16'd26155, 16'd19738};
                15'd9642 : data_rom <= {16'd26157, 16'd19736};
                15'd9643 : data_rom <= {16'd26159, 16'd19733};
                15'd9644 : data_rom <= {16'd26161, 16'd19731};
                15'd9645 : data_rom <= {16'd26163, 16'd19728};
                15'd9646 : data_rom <= {16'd26165, 16'd19726};
                15'd9647 : data_rom <= {16'd26167, 16'd19723};
                15'd9648 : data_rom <= {16'd26168, 16'd19721};
                15'd9649 : data_rom <= {16'd26170, 16'd19718};
                15'd9650 : data_rom <= {16'd26172, 16'd19716};
                15'd9651 : data_rom <= {16'd26174, 16'd19713};
                15'd9652 : data_rom <= {16'd26176, 16'd19711};
                15'd9653 : data_rom <= {16'd26178, 16'd19708};
                15'd9654 : data_rom <= {16'd26180, 16'd19706};
                15'd9655 : data_rom <= {16'd26182, 16'd19703};
                15'd9656 : data_rom <= {16'd26184, 16'd19701};
                15'd9657 : data_rom <= {16'd26186, 16'd19698};
                15'd9658 : data_rom <= {16'd26187, 16'd19696};
                15'd9659 : data_rom <= {16'd26189, 16'd19693};
                15'd9660 : data_rom <= {16'd26191, 16'd19691};
                15'd9661 : data_rom <= {16'd26193, 16'd19688};
                15'd9662 : data_rom <= {16'd26195, 16'd19686};
                15'd9663 : data_rom <= {16'd26197, 16'd19683};
                15'd9664 : data_rom <= {16'd26199, 16'd19681};
                15'd9665 : data_rom <= {16'd26201, 16'd19678};
                15'd9666 : data_rom <= {16'd26202, 16'd19675};
                15'd9667 : data_rom <= {16'd26204, 16'd19673};
                15'd9668 : data_rom <= {16'd26206, 16'd19670};
                15'd9669 : data_rom <= {16'd26208, 16'd19668};
                15'd9670 : data_rom <= {16'd26210, 16'd19665};
                15'd9671 : data_rom <= {16'd26212, 16'd19663};
                15'd9672 : data_rom <= {16'd26214, 16'd19660};
                15'd9673 : data_rom <= {16'd26216, 16'd19658};
                15'd9674 : data_rom <= {16'd26218, 16'd19655};
                15'd9675 : data_rom <= {16'd26219, 16'd19653};
                15'd9676 : data_rom <= {16'd26221, 16'd19650};
                15'd9677 : data_rom <= {16'd26223, 16'd19648};
                15'd9678 : data_rom <= {16'd26225, 16'd19645};
                15'd9679 : data_rom <= {16'd26227, 16'd19643};
                15'd9680 : data_rom <= {16'd26229, 16'd19640};
                15'd9681 : data_rom <= {16'd26231, 16'd19638};
                15'd9682 : data_rom <= {16'd26233, 16'd19635};
                15'd9683 : data_rom <= {16'd26235, 16'd19633};
                15'd9684 : data_rom <= {16'd26236, 16'd19630};
                15'd9685 : data_rom <= {16'd26238, 16'd19628};
                15'd9686 : data_rom <= {16'd26240, 16'd19625};
                15'd9687 : data_rom <= {16'd26242, 16'd19623};
                15'd9688 : data_rom <= {16'd26244, 16'd19620};
                15'd9689 : data_rom <= {16'd26246, 16'd19618};
                15'd9690 : data_rom <= {16'd26248, 16'd19615};
                15'd9691 : data_rom <= {16'd26250, 16'd19613};
                15'd9692 : data_rom <= {16'd26251, 16'd19610};
                15'd9693 : data_rom <= {16'd26253, 16'd19608};
                15'd9694 : data_rom <= {16'd26255, 16'd19605};
                15'd9695 : data_rom <= {16'd26257, 16'd19603};
                15'd9696 : data_rom <= {16'd26259, 16'd19600};
                15'd9697 : data_rom <= {16'd26261, 16'd19598};
                15'd9698 : data_rom <= {16'd26263, 16'd19595};
                15'd9699 : data_rom <= {16'd26265, 16'd19592};
                15'd9700 : data_rom <= {16'd26266, 16'd19590};
                15'd9701 : data_rom <= {16'd26268, 16'd19587};
                15'd9702 : data_rom <= {16'd26270, 16'd19585};
                15'd9703 : data_rom <= {16'd26272, 16'd19582};
                15'd9704 : data_rom <= {16'd26274, 16'd19580};
                15'd9705 : data_rom <= {16'd26276, 16'd19577};
                15'd9706 : data_rom <= {16'd26278, 16'd19575};
                15'd9707 : data_rom <= {16'd26280, 16'd19572};
                15'd9708 : data_rom <= {16'd26282, 16'd19570};
                15'd9709 : data_rom <= {16'd26283, 16'd19567};
                15'd9710 : data_rom <= {16'd26285, 16'd19565};
                15'd9711 : data_rom <= {16'd26287, 16'd19562};
                15'd9712 : data_rom <= {16'd26289, 16'd19560};
                15'd9713 : data_rom <= {16'd26291, 16'd19557};
                15'd9714 : data_rom <= {16'd26293, 16'd19555};
                15'd9715 : data_rom <= {16'd26295, 16'd19552};
                15'd9716 : data_rom <= {16'd26297, 16'd19550};
                15'd9717 : data_rom <= {16'd26298, 16'd19547};
                15'd9718 : data_rom <= {16'd26300, 16'd19545};
                15'd9719 : data_rom <= {16'd26302, 16'd19542};
                15'd9720 : data_rom <= {16'd26304, 16'd19540};
                15'd9721 : data_rom <= {16'd26306, 16'd19537};
                15'd9722 : data_rom <= {16'd26308, 16'd19535};
                15'd9723 : data_rom <= {16'd26310, 16'd19532};
                15'd9724 : data_rom <= {16'd26311, 16'd19529};
                15'd9725 : data_rom <= {16'd26313, 16'd19527};
                15'd9726 : data_rom <= {16'd26315, 16'd19524};
                15'd9727 : data_rom <= {16'd26317, 16'd19522};
                15'd9728 : data_rom <= {16'd26319, 16'd19519};
                15'd9729 : data_rom <= {16'd26321, 16'd19517};
                15'd9730 : data_rom <= {16'd26323, 16'd19514};
                15'd9731 : data_rom <= {16'd26325, 16'd19512};
                15'd9732 : data_rom <= {16'd26326, 16'd19509};
                15'd9733 : data_rom <= {16'd26328, 16'd19507};
                15'd9734 : data_rom <= {16'd26330, 16'd19504};
                15'd9735 : data_rom <= {16'd26332, 16'd19502};
                15'd9736 : data_rom <= {16'd26334, 16'd19499};
                15'd9737 : data_rom <= {16'd26336, 16'd19497};
                15'd9738 : data_rom <= {16'd26338, 16'd19494};
                15'd9739 : data_rom <= {16'd26340, 16'd19492};
                15'd9740 : data_rom <= {16'd26341, 16'd19489};
                15'd9741 : data_rom <= {16'd26343, 16'd19487};
                15'd9742 : data_rom <= {16'd26345, 16'd19484};
                15'd9743 : data_rom <= {16'd26347, 16'd19482};
                15'd9744 : data_rom <= {16'd26349, 16'd19479};
                15'd9745 : data_rom <= {16'd26351, 16'd19476};
                15'd9746 : data_rom <= {16'd26353, 16'd19474};
                15'd9747 : data_rom <= {16'd26355, 16'd19471};
                15'd9748 : data_rom <= {16'd26356, 16'd19469};
                15'd9749 : data_rom <= {16'd26358, 16'd19466};
                15'd9750 : data_rom <= {16'd26360, 16'd19464};
                15'd9751 : data_rom <= {16'd26362, 16'd19461};
                15'd9752 : data_rom <= {16'd26364, 16'd19459};
                15'd9753 : data_rom <= {16'd26366, 16'd19456};
                15'd9754 : data_rom <= {16'd26368, 16'd19454};
                15'd9755 : data_rom <= {16'd26369, 16'd19451};
                15'd9756 : data_rom <= {16'd26371, 16'd19449};
                15'd9757 : data_rom <= {16'd26373, 16'd19446};
                15'd9758 : data_rom <= {16'd26375, 16'd19444};
                15'd9759 : data_rom <= {16'd26377, 16'd19441};
                15'd9760 : data_rom <= {16'd26379, 16'd19439};
                15'd9761 : data_rom <= {16'd26381, 16'd19436};
                15'd9762 : data_rom <= {16'd26382, 16'd19434};
                15'd9763 : data_rom <= {16'd26384, 16'd19431};
                15'd9764 : data_rom <= {16'd26386, 16'd19428};
                15'd9765 : data_rom <= {16'd26388, 16'd19426};
                15'd9766 : data_rom <= {16'd26390, 16'd19423};
                15'd9767 : data_rom <= {16'd26392, 16'd19421};
                15'd9768 : data_rom <= {16'd26394, 16'd19418};
                15'd9769 : data_rom <= {16'd26396, 16'd19416};
                15'd9770 : data_rom <= {16'd26397, 16'd19413};
                15'd9771 : data_rom <= {16'd26399, 16'd19411};
                15'd9772 : data_rom <= {16'd26401, 16'd19408};
                15'd9773 : data_rom <= {16'd26403, 16'd19406};
                15'd9774 : data_rom <= {16'd26405, 16'd19403};
                15'd9775 : data_rom <= {16'd26407, 16'd19401};
                15'd9776 : data_rom <= {16'd26409, 16'd19398};
                15'd9777 : data_rom <= {16'd26410, 16'd19396};
                15'd9778 : data_rom <= {16'd26412, 16'd19393};
                15'd9779 : data_rom <= {16'd26414, 16'd19390};
                15'd9780 : data_rom <= {16'd26416, 16'd19388};
                15'd9781 : data_rom <= {16'd26418, 16'd19385};
                15'd9782 : data_rom <= {16'd26420, 16'd19383};
                15'd9783 : data_rom <= {16'd26422, 16'd19380};
                15'd9784 : data_rom <= {16'd26423, 16'd19378};
                15'd9785 : data_rom <= {16'd26425, 16'd19375};
                15'd9786 : data_rom <= {16'd26427, 16'd19373};
                15'd9787 : data_rom <= {16'd26429, 16'd19370};
                15'd9788 : data_rom <= {16'd26431, 16'd19368};
                15'd9789 : data_rom <= {16'd26433, 16'd19365};
                15'd9790 : data_rom <= {16'd26435, 16'd19363};
                15'd9791 : data_rom <= {16'd26436, 16'd19360};
                15'd9792 : data_rom <= {16'd26438, 16'd19358};
                15'd9793 : data_rom <= {16'd26440, 16'd19355};
                15'd9794 : data_rom <= {16'd26442, 16'd19352};
                15'd9795 : data_rom <= {16'd26444, 16'd19350};
                15'd9796 : data_rom <= {16'd26446, 16'd19347};
                15'd9797 : data_rom <= {16'd26448, 16'd19345};
                15'd9798 : data_rom <= {16'd26449, 16'd19342};
                15'd9799 : data_rom <= {16'd26451, 16'd19340};
                15'd9800 : data_rom <= {16'd26453, 16'd19337};
                15'd9801 : data_rom <= {16'd26455, 16'd19335};
                15'd9802 : data_rom <= {16'd26457, 16'd19332};
                15'd9803 : data_rom <= {16'd26459, 16'd19330};
                15'd9804 : data_rom <= {16'd26461, 16'd19327};
                15'd9805 : data_rom <= {16'd26462, 16'd19325};
                15'd9806 : data_rom <= {16'd26464, 16'd19322};
                15'd9807 : data_rom <= {16'd26466, 16'd19319};
                15'd9808 : data_rom <= {16'd26468, 16'd19317};
                15'd9809 : data_rom <= {16'd26470, 16'd19314};
                15'd9810 : data_rom <= {16'd26472, 16'd19312};
                15'd9811 : data_rom <= {16'd26473, 16'd19309};
                15'd9812 : data_rom <= {16'd26475, 16'd19307};
                15'd9813 : data_rom <= {16'd26477, 16'd19304};
                15'd9814 : data_rom <= {16'd26479, 16'd19302};
                15'd9815 : data_rom <= {16'd26481, 16'd19299};
                15'd9816 : data_rom <= {16'd26483, 16'd19297};
                15'd9817 : data_rom <= {16'd26485, 16'd19294};
                15'd9818 : data_rom <= {16'd26486, 16'd19292};
                15'd9819 : data_rom <= {16'd26488, 16'd19289};
                15'd9820 : data_rom <= {16'd26490, 16'd19286};
                15'd9821 : data_rom <= {16'd26492, 16'd19284};
                15'd9822 : data_rom <= {16'd26494, 16'd19281};
                15'd9823 : data_rom <= {16'd26496, 16'd19279};
                15'd9824 : data_rom <= {16'd26498, 16'd19276};
                15'd9825 : data_rom <= {16'd26499, 16'd19274};
                15'd9826 : data_rom <= {16'd26501, 16'd19271};
                15'd9827 : data_rom <= {16'd26503, 16'd19269};
                15'd9828 : data_rom <= {16'd26505, 16'd19266};
                15'd9829 : data_rom <= {16'd26507, 16'd19264};
                15'd9830 : data_rom <= {16'd26509, 16'd19261};
                15'd9831 : data_rom <= {16'd26510, 16'd19259};
                15'd9832 : data_rom <= {16'd26512, 16'd19256};
                15'd9833 : data_rom <= {16'd26514, 16'd19253};
                15'd9834 : data_rom <= {16'd26516, 16'd19251};
                15'd9835 : data_rom <= {16'd26518, 16'd19248};
                15'd9836 : data_rom <= {16'd26520, 16'd19246};
                15'd9837 : data_rom <= {16'd26522, 16'd19243};
                15'd9838 : data_rom <= {16'd26523, 16'd19241};
                15'd9839 : data_rom <= {16'd26525, 16'd19238};
                15'd9840 : data_rom <= {16'd26527, 16'd19236};
                15'd9841 : data_rom <= {16'd26529, 16'd19233};
                15'd9842 : data_rom <= {16'd26531, 16'd19231};
                15'd9843 : data_rom <= {16'd26533, 16'd19228};
                15'd9844 : data_rom <= {16'd26534, 16'd19225};
                15'd9845 : data_rom <= {16'd26536, 16'd19223};
                15'd9846 : data_rom <= {16'd26538, 16'd19220};
                15'd9847 : data_rom <= {16'd26540, 16'd19218};
                15'd9848 : data_rom <= {16'd26542, 16'd19215};
                15'd9849 : data_rom <= {16'd26544, 16'd19213};
                15'd9850 : data_rom <= {16'd26545, 16'd19210};
                15'd9851 : data_rom <= {16'd26547, 16'd19208};
                15'd9852 : data_rom <= {16'd26549, 16'd19205};
                15'd9853 : data_rom <= {16'd26551, 16'd19203};
                15'd9854 : data_rom <= {16'd26553, 16'd19200};
                15'd9855 : data_rom <= {16'd26555, 16'd19197};
                15'd9856 : data_rom <= {16'd26557, 16'd19195};
                15'd9857 : data_rom <= {16'd26558, 16'd19192};
                15'd9858 : data_rom <= {16'd26560, 16'd19190};
                15'd9859 : data_rom <= {16'd26562, 16'd19187};
                15'd9860 : data_rom <= {16'd26564, 16'd19185};
                15'd9861 : data_rom <= {16'd26566, 16'd19182};
                15'd9862 : data_rom <= {16'd26568, 16'd19180};
                15'd9863 : data_rom <= {16'd26569, 16'd19177};
                15'd9864 : data_rom <= {16'd26571, 16'd19175};
                15'd9865 : data_rom <= {16'd26573, 16'd19172};
                15'd9866 : data_rom <= {16'd26575, 16'd19169};
                15'd9867 : data_rom <= {16'd26577, 16'd19167};
                15'd9868 : data_rom <= {16'd26579, 16'd19164};
                15'd9869 : data_rom <= {16'd26580, 16'd19162};
                15'd9870 : data_rom <= {16'd26582, 16'd19159};
                15'd9871 : data_rom <= {16'd26584, 16'd19157};
                15'd9872 : data_rom <= {16'd26586, 16'd19154};
                15'd9873 : data_rom <= {16'd26588, 16'd19152};
                15'd9874 : data_rom <= {16'd26590, 16'd19149};
                15'd9875 : data_rom <= {16'd26591, 16'd19147};
                15'd9876 : data_rom <= {16'd26593, 16'd19144};
                15'd9877 : data_rom <= {16'd26595, 16'd19141};
                15'd9878 : data_rom <= {16'd26597, 16'd19139};
                15'd9879 : data_rom <= {16'd26599, 16'd19136};
                15'd9880 : data_rom <= {16'd26601, 16'd19134};
                15'd9881 : data_rom <= {16'd26602, 16'd19131};
                15'd9882 : data_rom <= {16'd26604, 16'd19129};
                15'd9883 : data_rom <= {16'd26606, 16'd19126};
                15'd9884 : data_rom <= {16'd26608, 16'd19124};
                15'd9885 : data_rom <= {16'd26610, 16'd19121};
                15'd9886 : data_rom <= {16'd26612, 16'd19118};
                15'd9887 : data_rom <= {16'd26613, 16'd19116};
                15'd9888 : data_rom <= {16'd26615, 16'd19113};
                15'd9889 : data_rom <= {16'd26617, 16'd19111};
                15'd9890 : data_rom <= {16'd26619, 16'd19108};
                15'd9891 : data_rom <= {16'd26621, 16'd19106};
                15'd9892 : data_rom <= {16'd26623, 16'd19103};
                15'd9893 : data_rom <= {16'd26624, 16'd19101};
                15'd9894 : data_rom <= {16'd26626, 16'd19098};
                15'd9895 : data_rom <= {16'd26628, 16'd19096};
                15'd9896 : data_rom <= {16'd26630, 16'd19093};
                15'd9897 : data_rom <= {16'd26632, 16'd19090};
                15'd9898 : data_rom <= {16'd26634, 16'd19088};
                15'd9899 : data_rom <= {16'd26635, 16'd19085};
                15'd9900 : data_rom <= {16'd26637, 16'd19083};
                15'd9901 : data_rom <= {16'd26639, 16'd19080};
                15'd9902 : data_rom <= {16'd26641, 16'd19078};
                15'd9903 : data_rom <= {16'd26643, 16'd19075};
                15'd9904 : data_rom <= {16'd26645, 16'd19073};
                15'd9905 : data_rom <= {16'd26646, 16'd19070};
                15'd9906 : data_rom <= {16'd26648, 16'd19067};
                15'd9907 : data_rom <= {16'd26650, 16'd19065};
                15'd9908 : data_rom <= {16'd26652, 16'd19062};
                15'd9909 : data_rom <= {16'd26654, 16'd19060};
                15'd9910 : data_rom <= {16'd26656, 16'd19057};
                15'd9911 : data_rom <= {16'd26657, 16'd19055};
                15'd9912 : data_rom <= {16'd26659, 16'd19052};
                15'd9913 : data_rom <= {16'd26661, 16'd19050};
                15'd9914 : data_rom <= {16'd26663, 16'd19047};
                15'd9915 : data_rom <= {16'd26665, 16'd19044};
                15'd9916 : data_rom <= {16'd26667, 16'd19042};
                15'd9917 : data_rom <= {16'd26668, 16'd19039};
                15'd9918 : data_rom <= {16'd26670, 16'd19037};
                15'd9919 : data_rom <= {16'd26672, 16'd19034};
                15'd9920 : data_rom <= {16'd26674, 16'd19032};
                15'd9921 : data_rom <= {16'd26676, 16'd19029};
                15'd9922 : data_rom <= {16'd26677, 16'd19027};
                15'd9923 : data_rom <= {16'd26679, 16'd19024};
                15'd9924 : data_rom <= {16'd26681, 16'd19021};
                15'd9925 : data_rom <= {16'd26683, 16'd19019};
                15'd9926 : data_rom <= {16'd26685, 16'd19016};
                15'd9927 : data_rom <= {16'd26687, 16'd19014};
                15'd9928 : data_rom <= {16'd26688, 16'd19011};
                15'd9929 : data_rom <= {16'd26690, 16'd19009};
                15'd9930 : data_rom <= {16'd26692, 16'd19006};
                15'd9931 : data_rom <= {16'd26694, 16'd19003};
                15'd9932 : data_rom <= {16'd26696, 16'd19001};
                15'd9933 : data_rom <= {16'd26698, 16'd18998};
                15'd9934 : data_rom <= {16'd26699, 16'd18996};
                15'd9935 : data_rom <= {16'd26701, 16'd18993};
                15'd9936 : data_rom <= {16'd26703, 16'd18991};
                15'd9937 : data_rom <= {16'd26705, 16'd18988};
                15'd9938 : data_rom <= {16'd26707, 16'd18986};
                15'd9939 : data_rom <= {16'd26708, 16'd18983};
                15'd9940 : data_rom <= {16'd26710, 16'd18980};
                15'd9941 : data_rom <= {16'd26712, 16'd18978};
                15'd9942 : data_rom <= {16'd26714, 16'd18975};
                15'd9943 : data_rom <= {16'd26716, 16'd18973};
                15'd9944 : data_rom <= {16'd26718, 16'd18970};
                15'd9945 : data_rom <= {16'd26719, 16'd18968};
                15'd9946 : data_rom <= {16'd26721, 16'd18965};
                15'd9947 : data_rom <= {16'd26723, 16'd18963};
                15'd9948 : data_rom <= {16'd26725, 16'd18960};
                15'd9949 : data_rom <= {16'd26727, 16'd18957};
                15'd9950 : data_rom <= {16'd26728, 16'd18955};
                15'd9951 : data_rom <= {16'd26730, 16'd18952};
                15'd9952 : data_rom <= {16'd26732, 16'd18950};
                15'd9953 : data_rom <= {16'd26734, 16'd18947};
                15'd9954 : data_rom <= {16'd26736, 16'd18945};
                15'd9955 : data_rom <= {16'd26738, 16'd18942};
                15'd9956 : data_rom <= {16'd26739, 16'd18939};
                15'd9957 : data_rom <= {16'd26741, 16'd18937};
                15'd9958 : data_rom <= {16'd26743, 16'd18934};
                15'd9959 : data_rom <= {16'd26745, 16'd18932};
                15'd9960 : data_rom <= {16'd26747, 16'd18929};
                15'd9961 : data_rom <= {16'd26748, 16'd18927};
                15'd9962 : data_rom <= {16'd26750, 16'd18924};
                15'd9963 : data_rom <= {16'd26752, 16'd18922};
                15'd9964 : data_rom <= {16'd26754, 16'd18919};
                15'd9965 : data_rom <= {16'd26756, 16'd18916};
                15'd9966 : data_rom <= {16'd26758, 16'd18914};
                15'd9967 : data_rom <= {16'd26759, 16'd18911};
                15'd9968 : data_rom <= {16'd26761, 16'd18909};
                15'd9969 : data_rom <= {16'd26763, 16'd18906};
                15'd9970 : data_rom <= {16'd26765, 16'd18904};
                15'd9971 : data_rom <= {16'd26767, 16'd18901};
                15'd9972 : data_rom <= {16'd26768, 16'd18898};
                15'd9973 : data_rom <= {16'd26770, 16'd18896};
                15'd9974 : data_rom <= {16'd26772, 16'd18893};
                15'd9975 : data_rom <= {16'd26774, 16'd18891};
                15'd9976 : data_rom <= {16'd26776, 16'd18888};
                15'd9977 : data_rom <= {16'd26777, 16'd18886};
                15'd9978 : data_rom <= {16'd26779, 16'd18883};
                15'd9979 : data_rom <= {16'd26781, 16'd18880};
                15'd9980 : data_rom <= {16'd26783, 16'd18878};
                15'd9981 : data_rom <= {16'd26785, 16'd18875};
                15'd9982 : data_rom <= {16'd26786, 16'd18873};
                15'd9983 : data_rom <= {16'd26788, 16'd18870};
                15'd9984 : data_rom <= {16'd26790, 16'd18868};
                15'd9985 : data_rom <= {16'd26792, 16'd18865};
                15'd9986 : data_rom <= {16'd26794, 16'd18862};
                15'd9987 : data_rom <= {16'd26796, 16'd18860};
                15'd9988 : data_rom <= {16'd26797, 16'd18857};
                15'd9989 : data_rom <= {16'd26799, 16'd18855};
                15'd9990 : data_rom <= {16'd26801, 16'd18852};
                15'd9991 : data_rom <= {16'd26803, 16'd18850};
                15'd9992 : data_rom <= {16'd26805, 16'd18847};
                15'd9993 : data_rom <= {16'd26806, 16'd18844};
                15'd9994 : data_rom <= {16'd26808, 16'd18842};
                15'd9995 : data_rom <= {16'd26810, 16'd18839};
                15'd9996 : data_rom <= {16'd26812, 16'd18837};
                15'd9997 : data_rom <= {16'd26814, 16'd18834};
                15'd9998 : data_rom <= {16'd26815, 16'd18832};
                15'd9999 : data_rom <= {16'd26817, 16'd18829};
                15'd10000 : data_rom <= {16'd26819, 16'd18826};
                15'd10001 : data_rom <= {16'd26821, 16'd18824};
                15'd10002 : data_rom <= {16'd26823, 16'd18821};
                15'd10003 : data_rom <= {16'd26824, 16'd18819};
                15'd10004 : data_rom <= {16'd26826, 16'd18816};
                15'd10005 : data_rom <= {16'd26828, 16'd18814};
                15'd10006 : data_rom <= {16'd26830, 16'd18811};
                15'd10007 : data_rom <= {16'd26832, 16'd18808};
                15'd10008 : data_rom <= {16'd26833, 16'd18806};
                15'd10009 : data_rom <= {16'd26835, 16'd18803};
                15'd10010 : data_rom <= {16'd26837, 16'd18801};
                15'd10011 : data_rom <= {16'd26839, 16'd18798};
                15'd10012 : data_rom <= {16'd26841, 16'd18796};
                15'd10013 : data_rom <= {16'd26842, 16'd18793};
                15'd10014 : data_rom <= {16'd26844, 16'd18790};
                15'd10015 : data_rom <= {16'd26846, 16'd18788};
                15'd10016 : data_rom <= {16'd26848, 16'd18785};
                15'd10017 : data_rom <= {16'd26850, 16'd18783};
                15'd10018 : data_rom <= {16'd26851, 16'd18780};
                15'd10019 : data_rom <= {16'd26853, 16'd18778};
                15'd10020 : data_rom <= {16'd26855, 16'd18775};
                15'd10021 : data_rom <= {16'd26857, 16'd18772};
                15'd10022 : data_rom <= {16'd26859, 16'd18770};
                15'd10023 : data_rom <= {16'd26860, 16'd18767};
                15'd10024 : data_rom <= {16'd26862, 16'd18765};
                15'd10025 : data_rom <= {16'd26864, 16'd18762};
                15'd10026 : data_rom <= {16'd26866, 16'd18760};
                15'd10027 : data_rom <= {16'd26868, 16'd18757};
                15'd10028 : data_rom <= {16'd26869, 16'd18754};
                15'd10029 : data_rom <= {16'd26871, 16'd18752};
                15'd10030 : data_rom <= {16'd26873, 16'd18749};
                15'd10031 : data_rom <= {16'd26875, 16'd18747};
                15'd10032 : data_rom <= {16'd26877, 16'd18744};
                15'd10033 : data_rom <= {16'd26878, 16'd18742};
                15'd10034 : data_rom <= {16'd26880, 16'd18739};
                15'd10035 : data_rom <= {16'd26882, 16'd18736};
                15'd10036 : data_rom <= {16'd26884, 16'd18734};
                15'd10037 : data_rom <= {16'd26886, 16'd18731};
                15'd10038 : data_rom <= {16'd26887, 16'd18729};
                15'd10039 : data_rom <= {16'd26889, 16'd18726};
                15'd10040 : data_rom <= {16'd26891, 16'd18723};
                15'd10041 : data_rom <= {16'd26893, 16'd18721};
                15'd10042 : data_rom <= {16'd26895, 16'd18718};
                15'd10043 : data_rom <= {16'd26896, 16'd18716};
                15'd10044 : data_rom <= {16'd26898, 16'd18713};
                15'd10045 : data_rom <= {16'd26900, 16'd18711};
                15'd10046 : data_rom <= {16'd26902, 16'd18708};
                15'd10047 : data_rom <= {16'd26904, 16'd18705};
                15'd10048 : data_rom <= {16'd26905, 16'd18703};
                15'd10049 : data_rom <= {16'd26907, 16'd18700};
                15'd10050 : data_rom <= {16'd26909, 16'd18698};
                15'd10051 : data_rom <= {16'd26911, 16'd18695};
                15'd10052 : data_rom <= {16'd26913, 16'd18693};
                15'd10053 : data_rom <= {16'd26914, 16'd18690};
                15'd10054 : data_rom <= {16'd26916, 16'd18687};
                15'd10055 : data_rom <= {16'd26918, 16'd18685};
                15'd10056 : data_rom <= {16'd26920, 16'd18682};
                15'd10057 : data_rom <= {16'd26921, 16'd18680};
                15'd10058 : data_rom <= {16'd26923, 16'd18677};
                15'd10059 : data_rom <= {16'd26925, 16'd18674};
                15'd10060 : data_rom <= {16'd26927, 16'd18672};
                15'd10061 : data_rom <= {16'd26929, 16'd18669};
                15'd10062 : data_rom <= {16'd26930, 16'd18667};
                15'd10063 : data_rom <= {16'd26932, 16'd18664};
                15'd10064 : data_rom <= {16'd26934, 16'd18662};
                15'd10065 : data_rom <= {16'd26936, 16'd18659};
                15'd10066 : data_rom <= {16'd26938, 16'd18656};
                15'd10067 : data_rom <= {16'd26939, 16'd18654};
                15'd10068 : data_rom <= {16'd26941, 16'd18651};
                15'd10069 : data_rom <= {16'd26943, 16'd18649};
                15'd10070 : data_rom <= {16'd26945, 16'd18646};
                15'd10071 : data_rom <= {16'd26947, 16'd18643};
                15'd10072 : data_rom <= {16'd26948, 16'd18641};
                15'd10073 : data_rom <= {16'd26950, 16'd18638};
                15'd10074 : data_rom <= {16'd26952, 16'd18636};
                15'd10075 : data_rom <= {16'd26954, 16'd18633};
                15'd10076 : data_rom <= {16'd26955, 16'd18631};
                15'd10077 : data_rom <= {16'd26957, 16'd18628};
                15'd10078 : data_rom <= {16'd26959, 16'd18625};
                15'd10079 : data_rom <= {16'd26961, 16'd18623};
                15'd10080 : data_rom <= {16'd26963, 16'd18620};
                15'd10081 : data_rom <= {16'd26964, 16'd18618};
                15'd10082 : data_rom <= {16'd26966, 16'd18615};
                15'd10083 : data_rom <= {16'd26968, 16'd18612};
                15'd10084 : data_rom <= {16'd26970, 16'd18610};
                15'd10085 : data_rom <= {16'd26972, 16'd18607};
                15'd10086 : data_rom <= {16'd26973, 16'd18605};
                15'd10087 : data_rom <= {16'd26975, 16'd18602};
                15'd10088 : data_rom <= {16'd26977, 16'd18600};
                15'd10089 : data_rom <= {16'd26979, 16'd18597};
                15'd10090 : data_rom <= {16'd26980, 16'd18594};
                15'd10091 : data_rom <= {16'd26982, 16'd18592};
                15'd10092 : data_rom <= {16'd26984, 16'd18589};
                15'd10093 : data_rom <= {16'd26986, 16'd18587};
                15'd10094 : data_rom <= {16'd26988, 16'd18584};
                15'd10095 : data_rom <= {16'd26989, 16'd18581};
                15'd10096 : data_rom <= {16'd26991, 16'd18579};
                15'd10097 : data_rom <= {16'd26993, 16'd18576};
                15'd10098 : data_rom <= {16'd26995, 16'd18574};
                15'd10099 : data_rom <= {16'd26996, 16'd18571};
                15'd10100 : data_rom <= {16'd26998, 16'd18568};
                15'd10101 : data_rom <= {16'd27000, 16'd18566};
                15'd10102 : data_rom <= {16'd27002, 16'd18563};
                15'd10103 : data_rom <= {16'd27004, 16'd18561};
                15'd10104 : data_rom <= {16'd27005, 16'd18558};
                15'd10105 : data_rom <= {16'd27007, 16'd18556};
                15'd10106 : data_rom <= {16'd27009, 16'd18553};
                15'd10107 : data_rom <= {16'd27011, 16'd18550};
                15'd10108 : data_rom <= {16'd27013, 16'd18548};
                15'd10109 : data_rom <= {16'd27014, 16'd18545};
                15'd10110 : data_rom <= {16'd27016, 16'd18543};
                15'd10111 : data_rom <= {16'd27018, 16'd18540};
                15'd10112 : data_rom <= {16'd27020, 16'd18537};
                15'd10113 : data_rom <= {16'd27021, 16'd18535};
                15'd10114 : data_rom <= {16'd27023, 16'd18532};
                15'd10115 : data_rom <= {16'd27025, 16'd18530};
                15'd10116 : data_rom <= {16'd27027, 16'd18527};
                15'd10117 : data_rom <= {16'd27029, 16'd18524};
                15'd10118 : data_rom <= {16'd27030, 16'd18522};
                15'd10119 : data_rom <= {16'd27032, 16'd18519};
                15'd10120 : data_rom <= {16'd27034, 16'd18517};
                15'd10121 : data_rom <= {16'd27036, 16'd18514};
                15'd10122 : data_rom <= {16'd27037, 16'd18512};
                15'd10123 : data_rom <= {16'd27039, 16'd18509};
                15'd10124 : data_rom <= {16'd27041, 16'd18506};
                15'd10125 : data_rom <= {16'd27043, 16'd18504};
                15'd10126 : data_rom <= {16'd27044, 16'd18501};
                15'd10127 : data_rom <= {16'd27046, 16'd18499};
                15'd10128 : data_rom <= {16'd27048, 16'd18496};
                15'd10129 : data_rom <= {16'd27050, 16'd18493};
                15'd10130 : data_rom <= {16'd27052, 16'd18491};
                15'd10131 : data_rom <= {16'd27053, 16'd18488};
                15'd10132 : data_rom <= {16'd27055, 16'd18486};
                15'd10133 : data_rom <= {16'd27057, 16'd18483};
                15'd10134 : data_rom <= {16'd27059, 16'd18480};
                15'd10135 : data_rom <= {16'd27060, 16'd18478};
                15'd10136 : data_rom <= {16'd27062, 16'd18475};
                15'd10137 : data_rom <= {16'd27064, 16'd18473};
                15'd10138 : data_rom <= {16'd27066, 16'd18470};
                15'd10139 : data_rom <= {16'd27068, 16'd18467};
                15'd10140 : data_rom <= {16'd27069, 16'd18465};
                15'd10141 : data_rom <= {16'd27071, 16'd18462};
                15'd10142 : data_rom <= {16'd27073, 16'd18460};
                15'd10143 : data_rom <= {16'd27075, 16'd18457};
                15'd10144 : data_rom <= {16'd27076, 16'd18454};
                15'd10145 : data_rom <= {16'd27078, 16'd18452};
                15'd10146 : data_rom <= {16'd27080, 16'd18449};
                15'd10147 : data_rom <= {16'd27082, 16'd18447};
                15'd10148 : data_rom <= {16'd27083, 16'd18444};
                15'd10149 : data_rom <= {16'd27085, 16'd18441};
                15'd10150 : data_rom <= {16'd27087, 16'd18439};
                15'd10151 : data_rom <= {16'd27089, 16'd18436};
                15'd10152 : data_rom <= {16'd27091, 16'd18434};
                15'd10153 : data_rom <= {16'd27092, 16'd18431};
                15'd10154 : data_rom <= {16'd27094, 16'd18428};
                15'd10155 : data_rom <= {16'd27096, 16'd18426};
                15'd10156 : data_rom <= {16'd27098, 16'd18423};
                15'd10157 : data_rom <= {16'd27099, 16'd18421};
                15'd10158 : data_rom <= {16'd27101, 16'd18418};
                15'd10159 : data_rom <= {16'd27103, 16'd18415};
                15'd10160 : data_rom <= {16'd27105, 16'd18413};
                15'd10161 : data_rom <= {16'd27106, 16'd18410};
                15'd10162 : data_rom <= {16'd27108, 16'd18408};
                15'd10163 : data_rom <= {16'd27110, 16'd18405};
                15'd10164 : data_rom <= {16'd27112, 16'd18402};
                15'd10165 : data_rom <= {16'd27113, 16'd18400};
                15'd10166 : data_rom <= {16'd27115, 16'd18397};
                15'd10167 : data_rom <= {16'd27117, 16'd18395};
                15'd10168 : data_rom <= {16'd27119, 16'd18392};
                15'd10169 : data_rom <= {16'd27121, 16'd18389};
                15'd10170 : data_rom <= {16'd27122, 16'd18387};
                15'd10171 : data_rom <= {16'd27124, 16'd18384};
                15'd10172 : data_rom <= {16'd27126, 16'd18382};
                15'd10173 : data_rom <= {16'd27128, 16'd18379};
                15'd10174 : data_rom <= {16'd27129, 16'd18376};
                15'd10175 : data_rom <= {16'd27131, 16'd18374};
                15'd10176 : data_rom <= {16'd27133, 16'd18371};
                15'd10177 : data_rom <= {16'd27135, 16'd18369};
                15'd10178 : data_rom <= {16'd27136, 16'd18366};
                15'd10179 : data_rom <= {16'd27138, 16'd18363};
                15'd10180 : data_rom <= {16'd27140, 16'd18361};
                15'd10181 : data_rom <= {16'd27142, 16'd18358};
                15'd10182 : data_rom <= {16'd27143, 16'd18356};
                15'd10183 : data_rom <= {16'd27145, 16'd18353};
                15'd10184 : data_rom <= {16'd27147, 16'd18350};
                15'd10185 : data_rom <= {16'd27149, 16'd18348};
                15'd10186 : data_rom <= {16'd27150, 16'd18345};
                15'd10187 : data_rom <= {16'd27152, 16'd18343};
                15'd10188 : data_rom <= {16'd27154, 16'd18340};
                15'd10189 : data_rom <= {16'd27156, 16'd18337};
                15'd10190 : data_rom <= {16'd27157, 16'd18335};
                15'd10191 : data_rom <= {16'd27159, 16'd18332};
                15'd10192 : data_rom <= {16'd27161, 16'd18330};
                15'd10193 : data_rom <= {16'd27163, 16'd18327};
                15'd10194 : data_rom <= {16'd27165, 16'd18324};
                15'd10195 : data_rom <= {16'd27166, 16'd18322};
                15'd10196 : data_rom <= {16'd27168, 16'd18319};
                15'd10197 : data_rom <= {16'd27170, 16'd18317};
                15'd10198 : data_rom <= {16'd27172, 16'd18314};
                15'd10199 : data_rom <= {16'd27173, 16'd18311};
                15'd10200 : data_rom <= {16'd27175, 16'd18309};
                15'd10201 : data_rom <= {16'd27177, 16'd18306};
                15'd10202 : data_rom <= {16'd27179, 16'd18304};
                15'd10203 : data_rom <= {16'd27180, 16'd18301};
                15'd10204 : data_rom <= {16'd27182, 16'd18298};
                15'd10205 : data_rom <= {16'd27184, 16'd18296};
                15'd10206 : data_rom <= {16'd27186, 16'd18293};
                15'd10207 : data_rom <= {16'd27187, 16'd18291};
                15'd10208 : data_rom <= {16'd27189, 16'd18288};
                15'd10209 : data_rom <= {16'd27191, 16'd18285};
                15'd10210 : data_rom <= {16'd27193, 16'd18283};
                15'd10211 : data_rom <= {16'd27194, 16'd18280};
                15'd10212 : data_rom <= {16'd27196, 16'd18278};
                15'd10213 : data_rom <= {16'd27198, 16'd18275};
                15'd10214 : data_rom <= {16'd27200, 16'd18272};
                15'd10215 : data_rom <= {16'd27201, 16'd18270};
                15'd10216 : data_rom <= {16'd27203, 16'd18267};
                15'd10217 : data_rom <= {16'd27205, 16'd18264};
                15'd10218 : data_rom <= {16'd27207, 16'd18262};
                15'd10219 : data_rom <= {16'd27208, 16'd18259};
                15'd10220 : data_rom <= {16'd27210, 16'd18257};
                15'd10221 : data_rom <= {16'd27212, 16'd18254};
                15'd10222 : data_rom <= {16'd27214, 16'd18251};
                15'd10223 : data_rom <= {16'd27215, 16'd18249};
                15'd10224 : data_rom <= {16'd27217, 16'd18246};
                15'd10225 : data_rom <= {16'd27219, 16'd18244};
                15'd10226 : data_rom <= {16'd27221, 16'd18241};
                15'd10227 : data_rom <= {16'd27222, 16'd18238};
                15'd10228 : data_rom <= {16'd27224, 16'd18236};
                15'd10229 : data_rom <= {16'd27226, 16'd18233};
                15'd10230 : data_rom <= {16'd27228, 16'd18231};
                15'd10231 : data_rom <= {16'd27229, 16'd18228};
                15'd10232 : data_rom <= {16'd27231, 16'd18225};
                15'd10233 : data_rom <= {16'd27233, 16'd18223};
                15'd10234 : data_rom <= {16'd27235, 16'd18220};
                15'd10235 : data_rom <= {16'd27236, 16'd18218};
                15'd10236 : data_rom <= {16'd27238, 16'd18215};
                15'd10237 : data_rom <= {16'd27240, 16'd18212};
                15'd10238 : data_rom <= {16'd27242, 16'd18210};
                15'd10239 : data_rom <= {16'd27243, 16'd18207};
                15'd10240 : data_rom <= {16'd27245, 16'd18204};
                15'd10241 : data_rom <= {16'd27247, 16'd18202};
                15'd10242 : data_rom <= {16'd27249, 16'd18199};
                15'd10243 : data_rom <= {16'd27250, 16'd18197};
                15'd10244 : data_rom <= {16'd27252, 16'd18194};
                15'd10245 : data_rom <= {16'd27254, 16'd18191};
                15'd10246 : data_rom <= {16'd27256, 16'd18189};
                15'd10247 : data_rom <= {16'd27257, 16'd18186};
                15'd10248 : data_rom <= {16'd27259, 16'd18184};
                15'd10249 : data_rom <= {16'd27261, 16'd18181};
                15'd10250 : data_rom <= {16'd27263, 16'd18178};
                15'd10251 : data_rom <= {16'd27264, 16'd18176};
                15'd10252 : data_rom <= {16'd27266, 16'd18173};
                15'd10253 : data_rom <= {16'd27268, 16'd18170};
                15'd10254 : data_rom <= {16'd27269, 16'd18168};
                15'd10255 : data_rom <= {16'd27271, 16'd18165};
                15'd10256 : data_rom <= {16'd27273, 16'd18163};
                15'd10257 : data_rom <= {16'd27275, 16'd18160};
                15'd10258 : data_rom <= {16'd27276, 16'd18157};
                15'd10259 : data_rom <= {16'd27278, 16'd18155};
                15'd10260 : data_rom <= {16'd27280, 16'd18152};
                15'd10261 : data_rom <= {16'd27282, 16'd18150};
                15'd10262 : data_rom <= {16'd27283, 16'd18147};
                15'd10263 : data_rom <= {16'd27285, 16'd18144};
                15'd10264 : data_rom <= {16'd27287, 16'd18142};
                15'd10265 : data_rom <= {16'd27289, 16'd18139};
                15'd10266 : data_rom <= {16'd27290, 16'd18136};
                15'd10267 : data_rom <= {16'd27292, 16'd18134};
                15'd10268 : data_rom <= {16'd27294, 16'd18131};
                15'd10269 : data_rom <= {16'd27296, 16'd18129};
                15'd10270 : data_rom <= {16'd27297, 16'd18126};
                15'd10271 : data_rom <= {16'd27299, 16'd18123};
                15'd10272 : data_rom <= {16'd27301, 16'd18121};
                15'd10273 : data_rom <= {16'd27303, 16'd18118};
                15'd10274 : data_rom <= {16'd27304, 16'd18116};
                15'd10275 : data_rom <= {16'd27306, 16'd18113};
                15'd10276 : data_rom <= {16'd27308, 16'd18110};
                15'd10277 : data_rom <= {16'd27309, 16'd18108};
                15'd10278 : data_rom <= {16'd27311, 16'd18105};
                15'd10279 : data_rom <= {16'd27313, 16'd18102};
                15'd10280 : data_rom <= {16'd27315, 16'd18100};
                15'd10281 : data_rom <= {16'd27316, 16'd18097};
                15'd10282 : data_rom <= {16'd27318, 16'd18095};
                15'd10283 : data_rom <= {16'd27320, 16'd18092};
                15'd10284 : data_rom <= {16'd27322, 16'd18089};
                15'd10285 : data_rom <= {16'd27323, 16'd18087};
                15'd10286 : data_rom <= {16'd27325, 16'd18084};
                15'd10287 : data_rom <= {16'd27327, 16'd18081};
                15'd10288 : data_rom <= {16'd27329, 16'd18079};
                15'd10289 : data_rom <= {16'd27330, 16'd18076};
                15'd10290 : data_rom <= {16'd27332, 16'd18074};
                15'd10291 : data_rom <= {16'd27334, 16'd18071};
                15'd10292 : data_rom <= {16'd27335, 16'd18068};
                15'd10293 : data_rom <= {16'd27337, 16'd18066};
                15'd10294 : data_rom <= {16'd27339, 16'd18063};
                15'd10295 : data_rom <= {16'd27341, 16'd18061};
                15'd10296 : data_rom <= {16'd27342, 16'd18058};
                15'd10297 : data_rom <= {16'd27344, 16'd18055};
                15'd10298 : data_rom <= {16'd27346, 16'd18053};
                15'd10299 : data_rom <= {16'd27348, 16'd18050};
                15'd10300 : data_rom <= {16'd27349, 16'd18047};
                15'd10301 : data_rom <= {16'd27351, 16'd18045};
                15'd10302 : data_rom <= {16'd27353, 16'd18042};
                15'd10303 : data_rom <= {16'd27355, 16'd18040};
                15'd10304 : data_rom <= {16'd27356, 16'd18037};
                15'd10305 : data_rom <= {16'd27358, 16'd18034};
                15'd10306 : data_rom <= {16'd27360, 16'd18032};
                15'd10307 : data_rom <= {16'd27361, 16'd18029};
                15'd10308 : data_rom <= {16'd27363, 16'd18026};
                15'd10309 : data_rom <= {16'd27365, 16'd18024};
                15'd10310 : data_rom <= {16'd27367, 16'd18021};
                15'd10311 : data_rom <= {16'd27368, 16'd18019};
                15'd10312 : data_rom <= {16'd27370, 16'd18016};
                15'd10313 : data_rom <= {16'd27372, 16'd18013};
                15'd10314 : data_rom <= {16'd27374, 16'd18011};
                15'd10315 : data_rom <= {16'd27375, 16'd18008};
                15'd10316 : data_rom <= {16'd27377, 16'd18005};
                15'd10317 : data_rom <= {16'd27379, 16'd18003};
                15'd10318 : data_rom <= {16'd27380, 16'd18000};
                15'd10319 : data_rom <= {16'd27382, 16'd17998};
                15'd10320 : data_rom <= {16'd27384, 16'd17995};
                15'd10321 : data_rom <= {16'd27386, 16'd17992};
                15'd10322 : data_rom <= {16'd27387, 16'd17990};
                15'd10323 : data_rom <= {16'd27389, 16'd17987};
                15'd10324 : data_rom <= {16'd27391, 16'd17984};
                15'd10325 : data_rom <= {16'd27393, 16'd17982};
                15'd10326 : data_rom <= {16'd27394, 16'd17979};
                15'd10327 : data_rom <= {16'd27396, 16'd17977};
                15'd10328 : data_rom <= {16'd27398, 16'd17974};
                15'd10329 : data_rom <= {16'd27399, 16'd17971};
                15'd10330 : data_rom <= {16'd27401, 16'd17969};
                15'd10331 : data_rom <= {16'd27403, 16'd17966};
                15'd10332 : data_rom <= {16'd27405, 16'd17963};
                15'd10333 : data_rom <= {16'd27406, 16'd17961};
                15'd10334 : data_rom <= {16'd27408, 16'd17958};
                15'd10335 : data_rom <= {16'd27410, 16'd17956};
                15'd10336 : data_rom <= {16'd27411, 16'd17953};
                15'd10337 : data_rom <= {16'd27413, 16'd17950};
                15'd10338 : data_rom <= {16'd27415, 16'd17948};
                15'd10339 : data_rom <= {16'd27417, 16'd17945};
                15'd10340 : data_rom <= {16'd27418, 16'd17942};
                15'd10341 : data_rom <= {16'd27420, 16'd17940};
                15'd10342 : data_rom <= {16'd27422, 16'd17937};
                15'd10343 : data_rom <= {16'd27424, 16'd17935};
                15'd10344 : data_rom <= {16'd27425, 16'd17932};
                15'd10345 : data_rom <= {16'd27427, 16'd17929};
                15'd10346 : data_rom <= {16'd27429, 16'd17927};
                15'd10347 : data_rom <= {16'd27430, 16'd17924};
                15'd10348 : data_rom <= {16'd27432, 16'd17921};
                15'd10349 : data_rom <= {16'd27434, 16'd17919};
                15'd10350 : data_rom <= {16'd27436, 16'd17916};
                15'd10351 : data_rom <= {16'd27437, 16'd17913};
                15'd10352 : data_rom <= {16'd27439, 16'd17911};
                15'd10353 : data_rom <= {16'd27441, 16'd17908};
                15'd10354 : data_rom <= {16'd27442, 16'd17906};
                15'd10355 : data_rom <= {16'd27444, 16'd17903};
                15'd10356 : data_rom <= {16'd27446, 16'd17900};
                15'd10357 : data_rom <= {16'd27448, 16'd17898};
                15'd10358 : data_rom <= {16'd27449, 16'd17895};
                15'd10359 : data_rom <= {16'd27451, 16'd17892};
                15'd10360 : data_rom <= {16'd27453, 16'd17890};
                15'd10361 : data_rom <= {16'd27454, 16'd17887};
                15'd10362 : data_rom <= {16'd27456, 16'd17885};
                15'd10363 : data_rom <= {16'd27458, 16'd17882};
                15'd10364 : data_rom <= {16'd27460, 16'd17879};
                15'd10365 : data_rom <= {16'd27461, 16'd17877};
                15'd10366 : data_rom <= {16'd27463, 16'd17874};
                15'd10367 : data_rom <= {16'd27465, 16'd17871};
                15'd10368 : data_rom <= {16'd27466, 16'd17869};
                15'd10369 : data_rom <= {16'd27468, 16'd17866};
                15'd10370 : data_rom <= {16'd27470, 16'd17863};
                15'd10371 : data_rom <= {16'd27472, 16'd17861};
                15'd10372 : data_rom <= {16'd27473, 16'd17858};
                15'd10373 : data_rom <= {16'd27475, 16'd17856};
                15'd10374 : data_rom <= {16'd27477, 16'd17853};
                15'd10375 : data_rom <= {16'd27478, 16'd17850};
                15'd10376 : data_rom <= {16'd27480, 16'd17848};
                15'd10377 : data_rom <= {16'd27482, 16'd17845};
                15'd10378 : data_rom <= {16'd27484, 16'd17842};
                15'd10379 : data_rom <= {16'd27485, 16'd17840};
                15'd10380 : data_rom <= {16'd27487, 16'd17837};
                15'd10381 : data_rom <= {16'd27489, 16'd17834};
                15'd10382 : data_rom <= {16'd27490, 16'd17832};
                15'd10383 : data_rom <= {16'd27492, 16'd17829};
                15'd10384 : data_rom <= {16'd27494, 16'd17827};
                15'd10385 : data_rom <= {16'd27496, 16'd17824};
                15'd10386 : data_rom <= {16'd27497, 16'd17821};
                15'd10387 : data_rom <= {16'd27499, 16'd17819};
                15'd10388 : data_rom <= {16'd27501, 16'd17816};
                15'd10389 : data_rom <= {16'd27502, 16'd17813};
                15'd10390 : data_rom <= {16'd27504, 16'd17811};
                15'd10391 : data_rom <= {16'd27506, 16'd17808};
                15'd10392 : data_rom <= {16'd27507, 16'd17805};
                15'd10393 : data_rom <= {16'd27509, 16'd17803};
                15'd10394 : data_rom <= {16'd27511, 16'd17800};
                15'd10395 : data_rom <= {16'd27513, 16'd17798};
                15'd10396 : data_rom <= {16'd27514, 16'd17795};
                15'd10397 : data_rom <= {16'd27516, 16'd17792};
                15'd10398 : data_rom <= {16'd27518, 16'd17790};
                15'd10399 : data_rom <= {16'd27519, 16'd17787};
                15'd10400 : data_rom <= {16'd27521, 16'd17784};
                15'd10401 : data_rom <= {16'd27523, 16'd17782};
                15'd10402 : data_rom <= {16'd27525, 16'd17779};
                15'd10403 : data_rom <= {16'd27526, 16'd17776};
                15'd10404 : data_rom <= {16'd27528, 16'd17774};
                15'd10405 : data_rom <= {16'd27530, 16'd17771};
                15'd10406 : data_rom <= {16'd27531, 16'd17769};
                15'd10407 : data_rom <= {16'd27533, 16'd17766};
                15'd10408 : data_rom <= {16'd27535, 16'd17763};
                15'd10409 : data_rom <= {16'd27536, 16'd17761};
                15'd10410 : data_rom <= {16'd27538, 16'd17758};
                15'd10411 : data_rom <= {16'd27540, 16'd17755};
                15'd10412 : data_rom <= {16'd27542, 16'd17753};
                15'd10413 : data_rom <= {16'd27543, 16'd17750};
                15'd10414 : data_rom <= {16'd27545, 16'd17747};
                15'd10415 : data_rom <= {16'd27547, 16'd17745};
                15'd10416 : data_rom <= {16'd27548, 16'd17742};
                15'd10417 : data_rom <= {16'd27550, 16'd17740};
                15'd10418 : data_rom <= {16'd27552, 16'd17737};
                15'd10419 : data_rom <= {16'd27553, 16'd17734};
                15'd10420 : data_rom <= {16'd27555, 16'd17732};
                15'd10421 : data_rom <= {16'd27557, 16'd17729};
                15'd10422 : data_rom <= {16'd27559, 16'd17726};
                15'd10423 : data_rom <= {16'd27560, 16'd17724};
                15'd10424 : data_rom <= {16'd27562, 16'd17721};
                15'd10425 : data_rom <= {16'd27564, 16'd17718};
                15'd10426 : data_rom <= {16'd27565, 16'd17716};
                15'd10427 : data_rom <= {16'd27567, 16'd17713};
                15'd10428 : data_rom <= {16'd27569, 16'd17710};
                15'd10429 : data_rom <= {16'd27570, 16'd17708};
                15'd10430 : data_rom <= {16'd27572, 16'd17705};
                15'd10431 : data_rom <= {16'd27574, 16'd17703};
                15'd10432 : data_rom <= {16'd27576, 16'd17700};
                15'd10433 : data_rom <= {16'd27577, 16'd17697};
                15'd10434 : data_rom <= {16'd27579, 16'd17695};
                15'd10435 : data_rom <= {16'd27581, 16'd17692};
                15'd10436 : data_rom <= {16'd27582, 16'd17689};
                15'd10437 : data_rom <= {16'd27584, 16'd17687};
                15'd10438 : data_rom <= {16'd27586, 16'd17684};
                15'd10439 : data_rom <= {16'd27587, 16'd17681};
                15'd10440 : data_rom <= {16'd27589, 16'd17679};
                15'd10441 : data_rom <= {16'd27591, 16'd17676};
                15'd10442 : data_rom <= {16'd27593, 16'd17673};
                15'd10443 : data_rom <= {16'd27594, 16'd17671};
                15'd10444 : data_rom <= {16'd27596, 16'd17668};
                15'd10445 : data_rom <= {16'd27598, 16'd17665};
                15'd10446 : data_rom <= {16'd27599, 16'd17663};
                15'd10447 : data_rom <= {16'd27601, 16'd17660};
                15'd10448 : data_rom <= {16'd27603, 16'd17658};
                15'd10449 : data_rom <= {16'd27604, 16'd17655};
                15'd10450 : data_rom <= {16'd27606, 16'd17652};
                15'd10451 : data_rom <= {16'd27608, 16'd17650};
                15'd10452 : data_rom <= {16'd27609, 16'd17647};
                15'd10453 : data_rom <= {16'd27611, 16'd17644};
                15'd10454 : data_rom <= {16'd27613, 16'd17642};
                15'd10455 : data_rom <= {16'd27615, 16'd17639};
                15'd10456 : data_rom <= {16'd27616, 16'd17636};
                15'd10457 : data_rom <= {16'd27618, 16'd17634};
                15'd10458 : data_rom <= {16'd27620, 16'd17631};
                15'd10459 : data_rom <= {16'd27621, 16'd17628};
                15'd10460 : data_rom <= {16'd27623, 16'd17626};
                15'd10461 : data_rom <= {16'd27625, 16'd17623};
                15'd10462 : data_rom <= {16'd27626, 16'd17620};
                15'd10463 : data_rom <= {16'd27628, 16'd17618};
                15'd10464 : data_rom <= {16'd27630, 16'd17615};
                15'd10465 : data_rom <= {16'd27631, 16'd17613};
                15'd10466 : data_rom <= {16'd27633, 16'd17610};
                15'd10467 : data_rom <= {16'd27635, 16'd17607};
                15'd10468 : data_rom <= {16'd27636, 16'd17605};
                15'd10469 : data_rom <= {16'd27638, 16'd17602};
                15'd10470 : data_rom <= {16'd27640, 16'd17599};
                15'd10471 : data_rom <= {16'd27642, 16'd17597};
                15'd10472 : data_rom <= {16'd27643, 16'd17594};
                15'd10473 : data_rom <= {16'd27645, 16'd17591};
                15'd10474 : data_rom <= {16'd27647, 16'd17589};
                15'd10475 : data_rom <= {16'd27648, 16'd17586};
                15'd10476 : data_rom <= {16'd27650, 16'd17583};
                15'd10477 : data_rom <= {16'd27652, 16'd17581};
                15'd10478 : data_rom <= {16'd27653, 16'd17578};
                15'd10479 : data_rom <= {16'd27655, 16'd17575};
                15'd10480 : data_rom <= {16'd27657, 16'd17573};
                15'd10481 : data_rom <= {16'd27658, 16'd17570};
                15'd10482 : data_rom <= {16'd27660, 16'd17567};
                15'd10483 : data_rom <= {16'd27662, 16'd17565};
                15'd10484 : data_rom <= {16'd27663, 16'd17562};
                15'd10485 : data_rom <= {16'd27665, 16'd17560};
                15'd10486 : data_rom <= {16'd27667, 16'd17557};
                15'd10487 : data_rom <= {16'd27669, 16'd17554};
                15'd10488 : data_rom <= {16'd27670, 16'd17552};
                15'd10489 : data_rom <= {16'd27672, 16'd17549};
                15'd10490 : data_rom <= {16'd27674, 16'd17546};
                15'd10491 : data_rom <= {16'd27675, 16'd17544};
                15'd10492 : data_rom <= {16'd27677, 16'd17541};
                15'd10493 : data_rom <= {16'd27679, 16'd17538};
                15'd10494 : data_rom <= {16'd27680, 16'd17536};
                15'd10495 : data_rom <= {16'd27682, 16'd17533};
                15'd10496 : data_rom <= {16'd27684, 16'd17530};
                15'd10497 : data_rom <= {16'd27685, 16'd17528};
                15'd10498 : data_rom <= {16'd27687, 16'd17525};
                15'd10499 : data_rom <= {16'd27689, 16'd17522};
                15'd10500 : data_rom <= {16'd27690, 16'd17520};
                15'd10501 : data_rom <= {16'd27692, 16'd17517};
                15'd10502 : data_rom <= {16'd27694, 16'd17514};
                15'd10503 : data_rom <= {16'd27695, 16'd17512};
                15'd10504 : data_rom <= {16'd27697, 16'd17509};
                15'd10505 : data_rom <= {16'd27699, 16'd17506};
                15'd10506 : data_rom <= {16'd27700, 16'd17504};
                15'd10507 : data_rom <= {16'd27702, 16'd17501};
                15'd10508 : data_rom <= {16'd27704, 16'd17498};
                15'd10509 : data_rom <= {16'd27705, 16'd17496};
                15'd10510 : data_rom <= {16'd27707, 16'd17493};
                15'd10511 : data_rom <= {16'd27709, 16'd17490};
                15'd10512 : data_rom <= {16'd27711, 16'd17488};
                15'd10513 : data_rom <= {16'd27712, 16'd17485};
                15'd10514 : data_rom <= {16'd27714, 16'd17483};
                15'd10515 : data_rom <= {16'd27716, 16'd17480};
                15'd10516 : data_rom <= {16'd27717, 16'd17477};
                15'd10517 : data_rom <= {16'd27719, 16'd17475};
                15'd10518 : data_rom <= {16'd27721, 16'd17472};
                15'd10519 : data_rom <= {16'd27722, 16'd17469};
                15'd10520 : data_rom <= {16'd27724, 16'd17467};
                15'd10521 : data_rom <= {16'd27726, 16'd17464};
                15'd10522 : data_rom <= {16'd27727, 16'd17461};
                15'd10523 : data_rom <= {16'd27729, 16'd17459};
                15'd10524 : data_rom <= {16'd27731, 16'd17456};
                15'd10525 : data_rom <= {16'd27732, 16'd17453};
                15'd10526 : data_rom <= {16'd27734, 16'd17451};
                15'd10527 : data_rom <= {16'd27736, 16'd17448};
                15'd10528 : data_rom <= {16'd27737, 16'd17445};
                15'd10529 : data_rom <= {16'd27739, 16'd17443};
                15'd10530 : data_rom <= {16'd27741, 16'd17440};
                15'd10531 : data_rom <= {16'd27742, 16'd17437};
                15'd10532 : data_rom <= {16'd27744, 16'd17435};
                15'd10533 : data_rom <= {16'd27746, 16'd17432};
                15'd10534 : data_rom <= {16'd27747, 16'd17429};
                15'd10535 : data_rom <= {16'd27749, 16'd17427};
                15'd10536 : data_rom <= {16'd27751, 16'd17424};
                15'd10537 : data_rom <= {16'd27752, 16'd17421};
                15'd10538 : data_rom <= {16'd27754, 16'd17419};
                15'd10539 : data_rom <= {16'd27756, 16'd17416};
                15'd10540 : data_rom <= {16'd27757, 16'd17413};
                15'd10541 : data_rom <= {16'd27759, 16'd17411};
                15'd10542 : data_rom <= {16'd27761, 16'd17408};
                15'd10543 : data_rom <= {16'd27762, 16'd17405};
                15'd10544 : data_rom <= {16'd27764, 16'd17403};
                15'd10545 : data_rom <= {16'd27766, 16'd17400};
                15'd10546 : data_rom <= {16'd27767, 16'd17397};
                15'd10547 : data_rom <= {16'd27769, 16'd17395};
                15'd10548 : data_rom <= {16'd27771, 16'd17392};
                15'd10549 : data_rom <= {16'd27772, 16'd17389};
                15'd10550 : data_rom <= {16'd27774, 16'd17387};
                15'd10551 : data_rom <= {16'd27776, 16'd17384};
                15'd10552 : data_rom <= {16'd27777, 16'd17381};
                15'd10553 : data_rom <= {16'd27779, 16'd17379};
                15'd10554 : data_rom <= {16'd27781, 16'd17376};
                15'd10555 : data_rom <= {16'd27782, 16'd17373};
                15'd10556 : data_rom <= {16'd27784, 16'd17371};
                15'd10557 : data_rom <= {16'd27786, 16'd17368};
                15'd10558 : data_rom <= {16'd27787, 16'd17365};
                15'd10559 : data_rom <= {16'd27789, 16'd17363};
                15'd10560 : data_rom <= {16'd27791, 16'd17360};
                15'd10561 : data_rom <= {16'd27792, 16'd17357};
                15'd10562 : data_rom <= {16'd27794, 16'd17355};
                15'd10563 : data_rom <= {16'd27796, 16'd17352};
                15'd10564 : data_rom <= {16'd27797, 16'd17349};
                15'd10565 : data_rom <= {16'd27799, 16'd17347};
                15'd10566 : data_rom <= {16'd27801, 16'd17344};
                15'd10567 : data_rom <= {16'd27802, 16'd17341};
                15'd10568 : data_rom <= {16'd27804, 16'd17339};
                15'd10569 : data_rom <= {16'd27806, 16'd17336};
                15'd10570 : data_rom <= {16'd27807, 16'd17333};
                15'd10571 : data_rom <= {16'd27809, 16'd17331};
                15'd10572 : data_rom <= {16'd27811, 16'd17328};
                15'd10573 : data_rom <= {16'd27812, 16'd17325};
                15'd10574 : data_rom <= {16'd27814, 16'd17323};
                15'd10575 : data_rom <= {16'd27816, 16'd17320};
                15'd10576 : data_rom <= {16'd27817, 16'd17317};
                15'd10577 : data_rom <= {16'd27819, 16'd17315};
                15'd10578 : data_rom <= {16'd27821, 16'd17312};
                15'd10579 : data_rom <= {16'd27822, 16'd17309};
                15'd10580 : data_rom <= {16'd27824, 16'd17307};
                15'd10581 : data_rom <= {16'd27826, 16'd17304};
                15'd10582 : data_rom <= {16'd27827, 16'd17301};
                15'd10583 : data_rom <= {16'd27829, 16'd17299};
                15'd10584 : data_rom <= {16'd27831, 16'd17296};
                15'd10585 : data_rom <= {16'd27832, 16'd17293};
                15'd10586 : data_rom <= {16'd27834, 16'd17291};
                15'd10587 : data_rom <= {16'd27836, 16'd17288};
                15'd10588 : data_rom <= {16'd27837, 16'd17285};
                15'd10589 : data_rom <= {16'd27839, 16'd17283};
                15'd10590 : data_rom <= {16'd27841, 16'd17280};
                15'd10591 : data_rom <= {16'd27842, 16'd17277};
                15'd10592 : data_rom <= {16'd27844, 16'd17275};
                15'd10593 : data_rom <= {16'd27845, 16'd17272};
                15'd10594 : data_rom <= {16'd27847, 16'd17269};
                15'd10595 : data_rom <= {16'd27849, 16'd17267};
                15'd10596 : data_rom <= {16'd27850, 16'd17264};
                15'd10597 : data_rom <= {16'd27852, 16'd17261};
                15'd10598 : data_rom <= {16'd27854, 16'd17259};
                15'd10599 : data_rom <= {16'd27855, 16'd17256};
                15'd10600 : data_rom <= {16'd27857, 16'd17253};
                15'd10601 : data_rom <= {16'd27859, 16'd17251};
                15'd10602 : data_rom <= {16'd27860, 16'd17248};
                15'd10603 : data_rom <= {16'd27862, 16'd17245};
                15'd10604 : data_rom <= {16'd27864, 16'd17243};
                15'd10605 : data_rom <= {16'd27865, 16'd17240};
                15'd10606 : data_rom <= {16'd27867, 16'd17237};
                15'd10607 : data_rom <= {16'd27869, 16'd17235};
                15'd10608 : data_rom <= {16'd27870, 16'd17232};
                15'd10609 : data_rom <= {16'd27872, 16'd17229};
                15'd10610 : data_rom <= {16'd27874, 16'd17227};
                15'd10611 : data_rom <= {16'd27875, 16'd17224};
                15'd10612 : data_rom <= {16'd27877, 16'd17221};
                15'd10613 : data_rom <= {16'd27879, 16'd17219};
                15'd10614 : data_rom <= {16'd27880, 16'd17216};
                15'd10615 : data_rom <= {16'd27882, 16'd17213};
                15'd10616 : data_rom <= {16'd27883, 16'd17211};
                15'd10617 : data_rom <= {16'd27885, 16'd17208};
                15'd10618 : data_rom <= {16'd27887, 16'd17205};
                15'd10619 : data_rom <= {16'd27888, 16'd17203};
                15'd10620 : data_rom <= {16'd27890, 16'd17200};
                15'd10621 : data_rom <= {16'd27892, 16'd17197};
                15'd10622 : data_rom <= {16'd27893, 16'd17195};
                15'd10623 : data_rom <= {16'd27895, 16'd17192};
                15'd10624 : data_rom <= {16'd27897, 16'd17189};
                15'd10625 : data_rom <= {16'd27898, 16'd17187};
                15'd10626 : data_rom <= {16'd27900, 16'd17184};
                15'd10627 : data_rom <= {16'd27902, 16'd17181};
                15'd10628 : data_rom <= {16'd27903, 16'd17179};
                15'd10629 : data_rom <= {16'd27905, 16'd17176};
                15'd10630 : data_rom <= {16'd27907, 16'd17173};
                15'd10631 : data_rom <= {16'd27908, 16'd17171};
                15'd10632 : data_rom <= {16'd27910, 16'd17168};
                15'd10633 : data_rom <= {16'd27912, 16'd17165};
                15'd10634 : data_rom <= {16'd27913, 16'd17163};
                15'd10635 : data_rom <= {16'd27915, 16'd17160};
                15'd10636 : data_rom <= {16'd27916, 16'd17157};
                15'd10637 : data_rom <= {16'd27918, 16'd17154};
                15'd10638 : data_rom <= {16'd27920, 16'd17152};
                15'd10639 : data_rom <= {16'd27921, 16'd17149};
                15'd10640 : data_rom <= {16'd27923, 16'd17146};
                15'd10641 : data_rom <= {16'd27925, 16'd17144};
                15'd10642 : data_rom <= {16'd27926, 16'd17141};
                15'd10643 : data_rom <= {16'd27928, 16'd17138};
                15'd10644 : data_rom <= {16'd27930, 16'd17136};
                15'd10645 : data_rom <= {16'd27931, 16'd17133};
                15'd10646 : data_rom <= {16'd27933, 16'd17130};
                15'd10647 : data_rom <= {16'd27935, 16'd17128};
                15'd10648 : data_rom <= {16'd27936, 16'd17125};
                15'd10649 : data_rom <= {16'd27938, 16'd17122};
                15'd10650 : data_rom <= {16'd27939, 16'd17120};
                15'd10651 : data_rom <= {16'd27941, 16'd17117};
                15'd10652 : data_rom <= {16'd27943, 16'd17114};
                15'd10653 : data_rom <= {16'd27944, 16'd17112};
                15'd10654 : data_rom <= {16'd27946, 16'd17109};
                15'd10655 : data_rom <= {16'd27948, 16'd17106};
                15'd10656 : data_rom <= {16'd27949, 16'd17104};
                15'd10657 : data_rom <= {16'd27951, 16'd17101};
                15'd10658 : data_rom <= {16'd27953, 16'd17098};
                15'd10659 : data_rom <= {16'd27954, 16'd17096};
                15'd10660 : data_rom <= {16'd27956, 16'd17093};
                15'd10661 : data_rom <= {16'd27957, 16'd17090};
                15'd10662 : data_rom <= {16'd27959, 16'd17088};
                15'd10663 : data_rom <= {16'd27961, 16'd17085};
                15'd10664 : data_rom <= {16'd27962, 16'd17082};
                15'd10665 : data_rom <= {16'd27964, 16'd17079};
                15'd10666 : data_rom <= {16'd27966, 16'd17077};
                15'd10667 : data_rom <= {16'd27967, 16'd17074};
                15'd10668 : data_rom <= {16'd27969, 16'd17071};
                15'd10669 : data_rom <= {16'd27971, 16'd17069};
                15'd10670 : data_rom <= {16'd27972, 16'd17066};
                15'd10671 : data_rom <= {16'd27974, 16'd17063};
                15'd10672 : data_rom <= {16'd27976, 16'd17061};
                15'd10673 : data_rom <= {16'd27977, 16'd17058};
                15'd10674 : data_rom <= {16'd27979, 16'd17055};
                15'd10675 : data_rom <= {16'd27980, 16'd17053};
                15'd10676 : data_rom <= {16'd27982, 16'd17050};
                15'd10677 : data_rom <= {16'd27984, 16'd17047};
                15'd10678 : data_rom <= {16'd27985, 16'd17045};
                15'd10679 : data_rom <= {16'd27987, 16'd17042};
                15'd10680 : data_rom <= {16'd27989, 16'd17039};
                15'd10681 : data_rom <= {16'd27990, 16'd17037};
                15'd10682 : data_rom <= {16'd27992, 16'd17034};
                15'd10683 : data_rom <= {16'd27993, 16'd17031};
                15'd10684 : data_rom <= {16'd27995, 16'd17029};
                15'd10685 : data_rom <= {16'd27997, 16'd17026};
                15'd10686 : data_rom <= {16'd27998, 16'd17023};
                15'd10687 : data_rom <= {16'd28000, 16'd17020};
                15'd10688 : data_rom <= {16'd28002, 16'd17018};
                15'd10689 : data_rom <= {16'd28003, 16'd17015};
                15'd10690 : data_rom <= {16'd28005, 16'd17012};
                15'd10691 : data_rom <= {16'd28007, 16'd17010};
                15'd10692 : data_rom <= {16'd28008, 16'd17007};
                15'd10693 : data_rom <= {16'd28010, 16'd17004};
                15'd10694 : data_rom <= {16'd28011, 16'd17002};
                15'd10695 : data_rom <= {16'd28013, 16'd16999};
                15'd10696 : data_rom <= {16'd28015, 16'd16996};
                15'd10697 : data_rom <= {16'd28016, 16'd16994};
                15'd10698 : data_rom <= {16'd28018, 16'd16991};
                15'd10699 : data_rom <= {16'd28020, 16'd16988};
                15'd10700 : data_rom <= {16'd28021, 16'd16986};
                15'd10701 : data_rom <= {16'd28023, 16'd16983};
                15'd10702 : data_rom <= {16'd28024, 16'd16980};
                15'd10703 : data_rom <= {16'd28026, 16'd16977};
                15'd10704 : data_rom <= {16'd28028, 16'd16975};
                15'd10705 : data_rom <= {16'd28029, 16'd16972};
                15'd10706 : data_rom <= {16'd28031, 16'd16969};
                15'd10707 : data_rom <= {16'd28033, 16'd16967};
                15'd10708 : data_rom <= {16'd28034, 16'd16964};
                15'd10709 : data_rom <= {16'd28036, 16'd16961};
                15'd10710 : data_rom <= {16'd28037, 16'd16959};
                15'd10711 : data_rom <= {16'd28039, 16'd16956};
                15'd10712 : data_rom <= {16'd28041, 16'd16953};
                15'd10713 : data_rom <= {16'd28042, 16'd16951};
                15'd10714 : data_rom <= {16'd28044, 16'd16948};
                15'd10715 : data_rom <= {16'd28046, 16'd16945};
                15'd10716 : data_rom <= {16'd28047, 16'd16943};
                15'd10717 : data_rom <= {16'd28049, 16'd16940};
                15'd10718 : data_rom <= {16'd28050, 16'd16937};
                15'd10719 : data_rom <= {16'd28052, 16'd16934};
                15'd10720 : data_rom <= {16'd28054, 16'd16932};
                15'd10721 : data_rom <= {16'd28055, 16'd16929};
                15'd10722 : data_rom <= {16'd28057, 16'd16926};
                15'd10723 : data_rom <= {16'd28059, 16'd16924};
                15'd10724 : data_rom <= {16'd28060, 16'd16921};
                15'd10725 : data_rom <= {16'd28062, 16'd16918};
                15'd10726 : data_rom <= {16'd28063, 16'd16916};
                15'd10727 : data_rom <= {16'd28065, 16'd16913};
                15'd10728 : data_rom <= {16'd28067, 16'd16910};
                15'd10729 : data_rom <= {16'd28068, 16'd16908};
                15'd10730 : data_rom <= {16'd28070, 16'd16905};
                15'd10731 : data_rom <= {16'd28072, 16'd16902};
                15'd10732 : data_rom <= {16'd28073, 16'd16900};
                15'd10733 : data_rom <= {16'd28075, 16'd16897};
                15'd10734 : data_rom <= {16'd28076, 16'd16894};
                15'd10735 : data_rom <= {16'd28078, 16'd16891};
                15'd10736 : data_rom <= {16'd28080, 16'd16889};
                15'd10737 : data_rom <= {16'd28081, 16'd16886};
                15'd10738 : data_rom <= {16'd28083, 16'd16883};
                15'd10739 : data_rom <= {16'd28085, 16'd16881};
                15'd10740 : data_rom <= {16'd28086, 16'd16878};
                15'd10741 : data_rom <= {16'd28088, 16'd16875};
                15'd10742 : data_rom <= {16'd28089, 16'd16873};
                15'd10743 : data_rom <= {16'd28091, 16'd16870};
                15'd10744 : data_rom <= {16'd28093, 16'd16867};
                15'd10745 : data_rom <= {16'd28094, 16'd16865};
                15'd10746 : data_rom <= {16'd28096, 16'd16862};
                15'd10747 : data_rom <= {16'd28097, 16'd16859};
                15'd10748 : data_rom <= {16'd28099, 16'd16856};
                15'd10749 : data_rom <= {16'd28101, 16'd16854};
                15'd10750 : data_rom <= {16'd28102, 16'd16851};
                15'd10751 : data_rom <= {16'd28104, 16'd16848};
                15'd10752 : data_rom <= {16'd28106, 16'd16846};
                15'd10753 : data_rom <= {16'd28107, 16'd16843};
                15'd10754 : data_rom <= {16'd28109, 16'd16840};
                15'd10755 : data_rom <= {16'd28110, 16'd16838};
                15'd10756 : data_rom <= {16'd28112, 16'd16835};
                15'd10757 : data_rom <= {16'd28114, 16'd16832};
                15'd10758 : data_rom <= {16'd28115, 16'd16829};
                15'd10759 : data_rom <= {16'd28117, 16'd16827};
                15'd10760 : data_rom <= {16'd28118, 16'd16824};
                15'd10761 : data_rom <= {16'd28120, 16'd16821};
                15'd10762 : data_rom <= {16'd28122, 16'd16819};
                15'd10763 : data_rom <= {16'd28123, 16'd16816};
                15'd10764 : data_rom <= {16'd28125, 16'd16813};
                15'd10765 : data_rom <= {16'd28127, 16'd16811};
                15'd10766 : data_rom <= {16'd28128, 16'd16808};
                15'd10767 : data_rom <= {16'd28130, 16'd16805};
                15'd10768 : data_rom <= {16'd28131, 16'd16803};
                15'd10769 : data_rom <= {16'd28133, 16'd16800};
                15'd10770 : data_rom <= {16'd28135, 16'd16797};
                15'd10771 : data_rom <= {16'd28136, 16'd16794};
                15'd10772 : data_rom <= {16'd28138, 16'd16792};
                15'd10773 : data_rom <= {16'd28139, 16'd16789};
                15'd10774 : data_rom <= {16'd28141, 16'd16786};
                15'd10775 : data_rom <= {16'd28143, 16'd16784};
                15'd10776 : data_rom <= {16'd28144, 16'd16781};
                15'd10777 : data_rom <= {16'd28146, 16'd16778};
                15'd10778 : data_rom <= {16'd28147, 16'd16776};
                15'd10779 : data_rom <= {16'd28149, 16'd16773};
                15'd10780 : data_rom <= {16'd28151, 16'd16770};
                15'd10781 : data_rom <= {16'd28152, 16'd16767};
                15'd10782 : data_rom <= {16'd28154, 16'd16765};
                15'd10783 : data_rom <= {16'd28155, 16'd16762};
                15'd10784 : data_rom <= {16'd28157, 16'd16759};
                15'd10785 : data_rom <= {16'd28159, 16'd16757};
                15'd10786 : data_rom <= {16'd28160, 16'd16754};
                15'd10787 : data_rom <= {16'd28162, 16'd16751};
                15'd10788 : data_rom <= {16'd28164, 16'd16749};
                15'd10789 : data_rom <= {16'd28165, 16'd16746};
                15'd10790 : data_rom <= {16'd28167, 16'd16743};
                15'd10791 : data_rom <= {16'd28168, 16'd16740};
                15'd10792 : data_rom <= {16'd28170, 16'd16738};
                15'd10793 : data_rom <= {16'd28172, 16'd16735};
                15'd10794 : data_rom <= {16'd28173, 16'd16732};
                15'd10795 : data_rom <= {16'd28175, 16'd16730};
                15'd10796 : data_rom <= {16'd28176, 16'd16727};
                15'd10797 : data_rom <= {16'd28178, 16'd16724};
                15'd10798 : data_rom <= {16'd28180, 16'd16722};
                15'd10799 : data_rom <= {16'd28181, 16'd16719};
                15'd10800 : data_rom <= {16'd28183, 16'd16716};
                15'd10801 : data_rom <= {16'd28184, 16'd16713};
                15'd10802 : data_rom <= {16'd28186, 16'd16711};
                15'd10803 : data_rom <= {16'd28188, 16'd16708};
                15'd10804 : data_rom <= {16'd28189, 16'd16705};
                15'd10805 : data_rom <= {16'd28191, 16'd16703};
                15'd10806 : data_rom <= {16'd28192, 16'd16700};
                15'd10807 : data_rom <= {16'd28194, 16'd16697};
                15'd10808 : data_rom <= {16'd28196, 16'd16695};
                15'd10809 : data_rom <= {16'd28197, 16'd16692};
                15'd10810 : data_rom <= {16'd28199, 16'd16689};
                15'd10811 : data_rom <= {16'd28200, 16'd16686};
                15'd10812 : data_rom <= {16'd28202, 16'd16684};
                15'd10813 : data_rom <= {16'd28204, 16'd16681};
                15'd10814 : data_rom <= {16'd28205, 16'd16678};
                15'd10815 : data_rom <= {16'd28207, 16'd16676};
                15'd10816 : data_rom <= {16'd28208, 16'd16673};
                15'd10817 : data_rom <= {16'd28210, 16'd16670};
                15'd10818 : data_rom <= {16'd28212, 16'd16667};
                15'd10819 : data_rom <= {16'd28213, 16'd16665};
                15'd10820 : data_rom <= {16'd28215, 16'd16662};
                15'd10821 : data_rom <= {16'd28216, 16'd16659};
                15'd10822 : data_rom <= {16'd28218, 16'd16657};
                15'd10823 : data_rom <= {16'd28220, 16'd16654};
                15'd10824 : data_rom <= {16'd28221, 16'd16651};
                15'd10825 : data_rom <= {16'd28223, 16'd16649};
                15'd10826 : data_rom <= {16'd28224, 16'd16646};
                15'd10827 : data_rom <= {16'd28226, 16'd16643};
                15'd10828 : data_rom <= {16'd28228, 16'd16640};
                15'd10829 : data_rom <= {16'd28229, 16'd16638};
                15'd10830 : data_rom <= {16'd28231, 16'd16635};
                15'd10831 : data_rom <= {16'd28232, 16'd16632};
                15'd10832 : data_rom <= {16'd28234, 16'd16630};
                15'd10833 : data_rom <= {16'd28236, 16'd16627};
                15'd10834 : data_rom <= {16'd28237, 16'd16624};
                15'd10835 : data_rom <= {16'd28239, 16'd16621};
                15'd10836 : data_rom <= {16'd28240, 16'd16619};
                15'd10837 : data_rom <= {16'd28242, 16'd16616};
                15'd10838 : data_rom <= {16'd28243, 16'd16613};
                15'd10839 : data_rom <= {16'd28245, 16'd16611};
                15'd10840 : data_rom <= {16'd28247, 16'd16608};
                15'd10841 : data_rom <= {16'd28248, 16'd16605};
                15'd10842 : data_rom <= {16'd28250, 16'd16603};
                15'd10843 : data_rom <= {16'd28251, 16'd16600};
                15'd10844 : data_rom <= {16'd28253, 16'd16597};
                15'd10845 : data_rom <= {16'd28255, 16'd16594};
                15'd10846 : data_rom <= {16'd28256, 16'd16592};
                15'd10847 : data_rom <= {16'd28258, 16'd16589};
                15'd10848 : data_rom <= {16'd28259, 16'd16586};
                15'd10849 : data_rom <= {16'd28261, 16'd16584};
                15'd10850 : data_rom <= {16'd28263, 16'd16581};
                15'd10851 : data_rom <= {16'd28264, 16'd16578};
                15'd10852 : data_rom <= {16'd28266, 16'd16575};
                15'd10853 : data_rom <= {16'd28267, 16'd16573};
                15'd10854 : data_rom <= {16'd28269, 16'd16570};
                15'd10855 : data_rom <= {16'd28271, 16'd16567};
                15'd10856 : data_rom <= {16'd28272, 16'd16565};
                15'd10857 : data_rom <= {16'd28274, 16'd16562};
                15'd10858 : data_rom <= {16'd28275, 16'd16559};
                15'd10859 : data_rom <= {16'd28277, 16'd16556};
                15'd10860 : data_rom <= {16'd28278, 16'd16554};
                15'd10861 : data_rom <= {16'd28280, 16'd16551};
                15'd10862 : data_rom <= {16'd28282, 16'd16548};
                15'd10863 : data_rom <= {16'd28283, 16'd16546};
                15'd10864 : data_rom <= {16'd28285, 16'd16543};
                15'd10865 : data_rom <= {16'd28286, 16'd16540};
                15'd10866 : data_rom <= {16'd28288, 16'd16537};
                15'd10867 : data_rom <= {16'd28290, 16'd16535};
                15'd10868 : data_rom <= {16'd28291, 16'd16532};
                15'd10869 : data_rom <= {16'd28293, 16'd16529};
                15'd10870 : data_rom <= {16'd28294, 16'd16527};
                15'd10871 : data_rom <= {16'd28296, 16'd16524};
                15'd10872 : data_rom <= {16'd28297, 16'd16521};
                15'd10873 : data_rom <= {16'd28299, 16'd16518};
                15'd10874 : data_rom <= {16'd28301, 16'd16516};
                15'd10875 : data_rom <= {16'd28302, 16'd16513};
                15'd10876 : data_rom <= {16'd28304, 16'd16510};
                15'd10877 : data_rom <= {16'd28305, 16'd16508};
                15'd10878 : data_rom <= {16'd28307, 16'd16505};
                15'd10879 : data_rom <= {16'd28309, 16'd16502};
                15'd10880 : data_rom <= {16'd28310, 16'd16499};
                15'd10881 : data_rom <= {16'd28312, 16'd16497};
                15'd10882 : data_rom <= {16'd28313, 16'd16494};
                15'd10883 : data_rom <= {16'd28315, 16'd16491};
                15'd10884 : data_rom <= {16'd28316, 16'd16489};
                15'd10885 : data_rom <= {16'd28318, 16'd16486};
                15'd10886 : data_rom <= {16'd28320, 16'd16483};
                15'd10887 : data_rom <= {16'd28321, 16'd16480};
                15'd10888 : data_rom <= {16'd28323, 16'd16478};
                15'd10889 : data_rom <= {16'd28324, 16'd16475};
                15'd10890 : data_rom <= {16'd28326, 16'd16472};
                15'd10891 : data_rom <= {16'd28328, 16'd16470};
                15'd10892 : data_rom <= {16'd28329, 16'd16467};
                15'd10893 : data_rom <= {16'd28331, 16'd16464};
                15'd10894 : data_rom <= {16'd28332, 16'd16461};
                15'd10895 : data_rom <= {16'd28334, 16'd16459};
                15'd10896 : data_rom <= {16'd28335, 16'd16456};
                15'd10897 : data_rom <= {16'd28337, 16'd16453};
                15'd10898 : data_rom <= {16'd28339, 16'd16451};
                15'd10899 : data_rom <= {16'd28340, 16'd16448};
                15'd10900 : data_rom <= {16'd28342, 16'd16445};
                15'd10901 : data_rom <= {16'd28343, 16'd16442};
                15'd10902 : data_rom <= {16'd28345, 16'd16440};
                15'd10903 : data_rom <= {16'd28346, 16'd16437};
                15'd10904 : data_rom <= {16'd28348, 16'd16434};
                15'd10905 : data_rom <= {16'd28350, 16'd16432};
                15'd10906 : data_rom <= {16'd28351, 16'd16429};
                15'd10907 : data_rom <= {16'd28353, 16'd16426};
                15'd10908 : data_rom <= {16'd28354, 16'd16423};
                15'd10909 : data_rom <= {16'd28356, 16'd16421};
                15'd10910 : data_rom <= {16'd28357, 16'd16418};
                15'd10911 : data_rom <= {16'd28359, 16'd16415};
                15'd10912 : data_rom <= {16'd28361, 16'd16413};
                15'd10913 : data_rom <= {16'd28362, 16'd16410};
                15'd10914 : data_rom <= {16'd28364, 16'd16407};
                15'd10915 : data_rom <= {16'd28365, 16'd16404};
                15'd10916 : data_rom <= {16'd28367, 16'd16402};
                15'd10917 : data_rom <= {16'd28368, 16'd16399};
                15'd10918 : data_rom <= {16'd28370, 16'd16396};
                15'd10919 : data_rom <= {16'd28372, 16'd16394};
                15'd10920 : data_rom <= {16'd28373, 16'd16391};
                15'd10921 : data_rom <= {16'd28375, 16'd16388};
                15'd10922 : data_rom <= {16'd28376, 16'd16385};
                15'd10923 : data_rom <= {16'd28378, 16'd16383};
                15'd10924 : data_rom <= {16'd28379, 16'd16380};
                15'd10925 : data_rom <= {16'd28381, 16'd16377};
                15'd10926 : data_rom <= {16'd28383, 16'd16374};
                15'd10927 : data_rom <= {16'd28384, 16'd16372};
                15'd10928 : data_rom <= {16'd28386, 16'd16369};
                15'd10929 : data_rom <= {16'd28387, 16'd16366};
                15'd10930 : data_rom <= {16'd28389, 16'd16364};
                15'd10931 : data_rom <= {16'd28390, 16'd16361};
                15'd10932 : data_rom <= {16'd28392, 16'd16358};
                15'd10933 : data_rom <= {16'd28394, 16'd16355};
                15'd10934 : data_rom <= {16'd28395, 16'd16353};
                15'd10935 : data_rom <= {16'd28397, 16'd16350};
                15'd10936 : data_rom <= {16'd28398, 16'd16347};
                15'd10937 : data_rom <= {16'd28400, 16'd16345};
                15'd10938 : data_rom <= {16'd28401, 16'd16342};
                15'd10939 : data_rom <= {16'd28403, 16'd16339};
                15'd10940 : data_rom <= {16'd28405, 16'd16336};
                15'd10941 : data_rom <= {16'd28406, 16'd16334};
                15'd10942 : data_rom <= {16'd28408, 16'd16331};
                15'd10943 : data_rom <= {16'd28409, 16'd16328};
                15'd10944 : data_rom <= {16'd28411, 16'd16325};
                15'd10945 : data_rom <= {16'd28412, 16'd16323};
                15'd10946 : data_rom <= {16'd28414, 16'd16320};
                15'd10947 : data_rom <= {16'd28416, 16'd16317};
                15'd10948 : data_rom <= {16'd28417, 16'd16315};
                15'd10949 : data_rom <= {16'd28419, 16'd16312};
                15'd10950 : data_rom <= {16'd28420, 16'd16309};
                15'd10951 : data_rom <= {16'd28422, 16'd16306};
                15'd10952 : data_rom <= {16'd28423, 16'd16304};
                15'd10953 : data_rom <= {16'd28425, 16'd16301};
                15'd10954 : data_rom <= {16'd28426, 16'd16298};
                15'd10955 : data_rom <= {16'd28428, 16'd16295};
                15'd10956 : data_rom <= {16'd28430, 16'd16293};
                15'd10957 : data_rom <= {16'd28431, 16'd16290};
                15'd10958 : data_rom <= {16'd28433, 16'd16287};
                15'd10959 : data_rom <= {16'd28434, 16'd16285};
                15'd10960 : data_rom <= {16'd28436, 16'd16282};
                15'd10961 : data_rom <= {16'd28437, 16'd16279};
                15'd10962 : data_rom <= {16'd28439, 16'd16276};
                15'd10963 : data_rom <= {16'd28441, 16'd16274};
                15'd10964 : data_rom <= {16'd28442, 16'd16271};
                15'd10965 : data_rom <= {16'd28444, 16'd16268};
                15'd10966 : data_rom <= {16'd28445, 16'd16265};
                15'd10967 : data_rom <= {16'd28447, 16'd16263};
                15'd10968 : data_rom <= {16'd28448, 16'd16260};
                15'd10969 : data_rom <= {16'd28450, 16'd16257};
                15'd10970 : data_rom <= {16'd28451, 16'd16255};
                15'd10971 : data_rom <= {16'd28453, 16'd16252};
                15'd10972 : data_rom <= {16'd28455, 16'd16249};
                15'd10973 : data_rom <= {16'd28456, 16'd16246};
                15'd10974 : data_rom <= {16'd28458, 16'd16244};
                15'd10975 : data_rom <= {16'd28459, 16'd16241};
                15'd10976 : data_rom <= {16'd28461, 16'd16238};
                15'd10977 : data_rom <= {16'd28462, 16'd16235};
                15'd10978 : data_rom <= {16'd28464, 16'd16233};
                15'd10979 : data_rom <= {16'd28465, 16'd16230};
                15'd10980 : data_rom <= {16'd28467, 16'd16227};
                15'd10981 : data_rom <= {16'd28469, 16'd16225};
                15'd10982 : data_rom <= {16'd28470, 16'd16222};
                15'd10983 : data_rom <= {16'd28472, 16'd16219};
                15'd10984 : data_rom <= {16'd28473, 16'd16216};
                15'd10985 : data_rom <= {16'd28475, 16'd16214};
                15'd10986 : data_rom <= {16'd28476, 16'd16211};
                15'd10987 : data_rom <= {16'd28478, 16'd16208};
                15'd10988 : data_rom <= {16'd28479, 16'd16205};
                15'd10989 : data_rom <= {16'd28481, 16'd16203};
                15'd10990 : data_rom <= {16'd28483, 16'd16200};
                15'd10991 : data_rom <= {16'd28484, 16'd16197};
                15'd10992 : data_rom <= {16'd28486, 16'd16195};
                15'd10993 : data_rom <= {16'd28487, 16'd16192};
                15'd10994 : data_rom <= {16'd28489, 16'd16189};
                15'd10995 : data_rom <= {16'd28490, 16'd16186};
                15'd10996 : data_rom <= {16'd28492, 16'd16184};
                15'd10997 : data_rom <= {16'd28493, 16'd16181};
                15'd10998 : data_rom <= {16'd28495, 16'd16178};
                15'd10999 : data_rom <= {16'd28497, 16'd16175};
                15'd11000 : data_rom <= {16'd28498, 16'd16173};
                15'd11001 : data_rom <= {16'd28500, 16'd16170};
                15'd11002 : data_rom <= {16'd28501, 16'd16167};
                15'd11003 : data_rom <= {16'd28503, 16'd16164};
                15'd11004 : data_rom <= {16'd28504, 16'd16162};
                15'd11005 : data_rom <= {16'd28506, 16'd16159};
                15'd11006 : data_rom <= {16'd28507, 16'd16156};
                15'd11007 : data_rom <= {16'd28509, 16'd16154};
                15'd11008 : data_rom <= {16'd28510, 16'd16151};
                15'd11009 : data_rom <= {16'd28512, 16'd16148};
                15'd11010 : data_rom <= {16'd28514, 16'd16145};
                15'd11011 : data_rom <= {16'd28515, 16'd16143};
                15'd11012 : data_rom <= {16'd28517, 16'd16140};
                15'd11013 : data_rom <= {16'd28518, 16'd16137};
                15'd11014 : data_rom <= {16'd28520, 16'd16134};
                15'd11015 : data_rom <= {16'd28521, 16'd16132};
                15'd11016 : data_rom <= {16'd28523, 16'd16129};
                15'd11017 : data_rom <= {16'd28524, 16'd16126};
                15'd11018 : data_rom <= {16'd28526, 16'd16123};
                15'd11019 : data_rom <= {16'd28528, 16'd16121};
                15'd11020 : data_rom <= {16'd28529, 16'd16118};
                15'd11021 : data_rom <= {16'd28531, 16'd16115};
                15'd11022 : data_rom <= {16'd28532, 16'd16113};
                15'd11023 : data_rom <= {16'd28534, 16'd16110};
                15'd11024 : data_rom <= {16'd28535, 16'd16107};
                15'd11025 : data_rom <= {16'd28537, 16'd16104};
                15'd11026 : data_rom <= {16'd28538, 16'd16102};
                15'd11027 : data_rom <= {16'd28540, 16'd16099};
                15'd11028 : data_rom <= {16'd28541, 16'd16096};
                15'd11029 : data_rom <= {16'd28543, 16'd16093};
                15'd11030 : data_rom <= {16'd28544, 16'd16091};
                15'd11031 : data_rom <= {16'd28546, 16'd16088};
                15'd11032 : data_rom <= {16'd28548, 16'd16085};
                15'd11033 : data_rom <= {16'd28549, 16'd16082};
                15'd11034 : data_rom <= {16'd28551, 16'd16080};
                15'd11035 : data_rom <= {16'd28552, 16'd16077};
                15'd11036 : data_rom <= {16'd28554, 16'd16074};
                15'd11037 : data_rom <= {16'd28555, 16'd16071};
                15'd11038 : data_rom <= {16'd28557, 16'd16069};
                15'd11039 : data_rom <= {16'd28558, 16'd16066};
                15'd11040 : data_rom <= {16'd28560, 16'd16063};
                15'd11041 : data_rom <= {16'd28561, 16'd16061};
                15'd11042 : data_rom <= {16'd28563, 16'd16058};
                15'd11043 : data_rom <= {16'd28565, 16'd16055};
                15'd11044 : data_rom <= {16'd28566, 16'd16052};
                15'd11045 : data_rom <= {16'd28568, 16'd16050};
                15'd11046 : data_rom <= {16'd28569, 16'd16047};
                15'd11047 : data_rom <= {16'd28571, 16'd16044};
                15'd11048 : data_rom <= {16'd28572, 16'd16041};
                15'd11049 : data_rom <= {16'd28574, 16'd16039};
                15'd11050 : data_rom <= {16'd28575, 16'd16036};
                15'd11051 : data_rom <= {16'd28577, 16'd16033};
                15'd11052 : data_rom <= {16'd28578, 16'd16030};
                15'd11053 : data_rom <= {16'd28580, 16'd16028};
                15'd11054 : data_rom <= {16'd28581, 16'd16025};
                15'd11055 : data_rom <= {16'd28583, 16'd16022};
                15'd11056 : data_rom <= {16'd28585, 16'd16019};
                15'd11057 : data_rom <= {16'd28586, 16'd16017};
                15'd11058 : data_rom <= {16'd28588, 16'd16014};
                15'd11059 : data_rom <= {16'd28589, 16'd16011};
                15'd11060 : data_rom <= {16'd28591, 16'd16008};
                15'd11061 : data_rom <= {16'd28592, 16'd16006};
                15'd11062 : data_rom <= {16'd28594, 16'd16003};
                15'd11063 : data_rom <= {16'd28595, 16'd16000};
                15'd11064 : data_rom <= {16'd28597, 16'd15998};
                15'd11065 : data_rom <= {16'd28598, 16'd15995};
                15'd11066 : data_rom <= {16'd28600, 16'd15992};
                15'd11067 : data_rom <= {16'd28601, 16'd15989};
                15'd11068 : data_rom <= {16'd28603, 16'd15987};
                15'd11069 : data_rom <= {16'd28604, 16'd15984};
                15'd11070 : data_rom <= {16'd28606, 16'd15981};
                15'd11071 : data_rom <= {16'd28608, 16'd15978};
                15'd11072 : data_rom <= {16'd28609, 16'd15976};
                15'd11073 : data_rom <= {16'd28611, 16'd15973};
                15'd11074 : data_rom <= {16'd28612, 16'd15970};
                15'd11075 : data_rom <= {16'd28614, 16'd15967};
                15'd11076 : data_rom <= {16'd28615, 16'd15965};
                15'd11077 : data_rom <= {16'd28617, 16'd15962};
                15'd11078 : data_rom <= {16'd28618, 16'd15959};
                15'd11079 : data_rom <= {16'd28620, 16'd15956};
                15'd11080 : data_rom <= {16'd28621, 16'd15954};
                15'd11081 : data_rom <= {16'd28623, 16'd15951};
                15'd11082 : data_rom <= {16'd28624, 16'd15948};
                15'd11083 : data_rom <= {16'd28626, 16'd15945};
                15'd11084 : data_rom <= {16'd28627, 16'd15943};
                15'd11085 : data_rom <= {16'd28629, 16'd15940};
                15'd11086 : data_rom <= {16'd28630, 16'd15937};
                15'd11087 : data_rom <= {16'd28632, 16'd15934};
                15'd11088 : data_rom <= {16'd28634, 16'd15932};
                15'd11089 : data_rom <= {16'd28635, 16'd15929};
                15'd11090 : data_rom <= {16'd28637, 16'd15926};
                15'd11091 : data_rom <= {16'd28638, 16'd15923};
                15'd11092 : data_rom <= {16'd28640, 16'd15921};
                15'd11093 : data_rom <= {16'd28641, 16'd15918};
                15'd11094 : data_rom <= {16'd28643, 16'd15915};
                15'd11095 : data_rom <= {16'd28644, 16'd15912};
                15'd11096 : data_rom <= {16'd28646, 16'd15910};
                15'd11097 : data_rom <= {16'd28647, 16'd15907};
                15'd11098 : data_rom <= {16'd28649, 16'd15904};
                15'd11099 : data_rom <= {16'd28650, 16'd15901};
                15'd11100 : data_rom <= {16'd28652, 16'd15899};
                15'd11101 : data_rom <= {16'd28653, 16'd15896};
                15'd11102 : data_rom <= {16'd28655, 16'd15893};
                15'd11103 : data_rom <= {16'd28656, 16'd15890};
                15'd11104 : data_rom <= {16'd28658, 16'd15888};
                15'd11105 : data_rom <= {16'd28659, 16'd15885};
                15'd11106 : data_rom <= {16'd28661, 16'd15882};
                15'd11107 : data_rom <= {16'd28663, 16'd15879};
                15'd11108 : data_rom <= {16'd28664, 16'd15877};
                15'd11109 : data_rom <= {16'd28666, 16'd15874};
                15'd11110 : data_rom <= {16'd28667, 16'd15871};
                15'd11111 : data_rom <= {16'd28669, 16'd15868};
                15'd11112 : data_rom <= {16'd28670, 16'd15866};
                15'd11113 : data_rom <= {16'd28672, 16'd15863};
                15'd11114 : data_rom <= {16'd28673, 16'd15860};
                15'd11115 : data_rom <= {16'd28675, 16'd15857};
                15'd11116 : data_rom <= {16'd28676, 16'd15855};
                15'd11117 : data_rom <= {16'd28678, 16'd15852};
                15'd11118 : data_rom <= {16'd28679, 16'd15849};
                15'd11119 : data_rom <= {16'd28681, 16'd15846};
                15'd11120 : data_rom <= {16'd28682, 16'd15844};
                15'd11121 : data_rom <= {16'd28684, 16'd15841};
                15'd11122 : data_rom <= {16'd28685, 16'd15838};
                15'd11123 : data_rom <= {16'd28687, 16'd15835};
                15'd11124 : data_rom <= {16'd28688, 16'd15833};
                15'd11125 : data_rom <= {16'd28690, 16'd15830};
                15'd11126 : data_rom <= {16'd28691, 16'd15827};
                15'd11127 : data_rom <= {16'd28693, 16'd15824};
                15'd11128 : data_rom <= {16'd28694, 16'd15822};
                15'd11129 : data_rom <= {16'd28696, 16'd15819};
                15'd11130 : data_rom <= {16'd28697, 16'd15816};
                15'd11131 : data_rom <= {16'd28699, 16'd15813};
                15'd11132 : data_rom <= {16'd28700, 16'd15811};
                15'd11133 : data_rom <= {16'd28702, 16'd15808};
                15'd11134 : data_rom <= {16'd28704, 16'd15805};
                15'd11135 : data_rom <= {16'd28705, 16'd15802};
                15'd11136 : data_rom <= {16'd28707, 16'd15800};
                15'd11137 : data_rom <= {16'd28708, 16'd15797};
                15'd11138 : data_rom <= {16'd28710, 16'd15794};
                15'd11139 : data_rom <= {16'd28711, 16'd15791};
                15'd11140 : data_rom <= {16'd28713, 16'd15789};
                15'd11141 : data_rom <= {16'd28714, 16'd15786};
                15'd11142 : data_rom <= {16'd28716, 16'd15783};
                15'd11143 : data_rom <= {16'd28717, 16'd15780};
                15'd11144 : data_rom <= {16'd28719, 16'd15778};
                15'd11145 : data_rom <= {16'd28720, 16'd15775};
                15'd11146 : data_rom <= {16'd28722, 16'd15772};
                15'd11147 : data_rom <= {16'd28723, 16'd15769};
                15'd11148 : data_rom <= {16'd28725, 16'd15767};
                15'd11149 : data_rom <= {16'd28726, 16'd15764};
                15'd11150 : data_rom <= {16'd28728, 16'd15761};
                15'd11151 : data_rom <= {16'd28729, 16'd15758};
                15'd11152 : data_rom <= {16'd28731, 16'd15756};
                15'd11153 : data_rom <= {16'd28732, 16'd15753};
                15'd11154 : data_rom <= {16'd28734, 16'd15750};
                15'd11155 : data_rom <= {16'd28735, 16'd15747};
                15'd11156 : data_rom <= {16'd28737, 16'd15745};
                15'd11157 : data_rom <= {16'd28738, 16'd15742};
                15'd11158 : data_rom <= {16'd28740, 16'd15739};
                15'd11159 : data_rom <= {16'd28741, 16'd15736};
                15'd11160 : data_rom <= {16'd28743, 16'd15734};
                15'd11161 : data_rom <= {16'd28744, 16'd15731};
                15'd11162 : data_rom <= {16'd28746, 16'd15728};
                15'd11163 : data_rom <= {16'd28747, 16'd15725};
                15'd11164 : data_rom <= {16'd28749, 16'd15723};
                15'd11165 : data_rom <= {16'd28750, 16'd15720};
                15'd11166 : data_rom <= {16'd28752, 16'd15717};
                15'd11167 : data_rom <= {16'd28753, 16'd15714};
                15'd11168 : data_rom <= {16'd28755, 16'd15712};
                15'd11169 : data_rom <= {16'd28756, 16'd15709};
                15'd11170 : data_rom <= {16'd28758, 16'd15706};
                15'd11171 : data_rom <= {16'd28759, 16'd15703};
                15'd11172 : data_rom <= {16'd28761, 16'd15701};
                15'd11173 : data_rom <= {16'd28762, 16'd15698};
                15'd11174 : data_rom <= {16'd28764, 16'd15695};
                15'd11175 : data_rom <= {16'd28765, 16'd15692};
                15'd11176 : data_rom <= {16'd28767, 16'd15690};
                15'd11177 : data_rom <= {16'd28768, 16'd15687};
                15'd11178 : data_rom <= {16'd28770, 16'd15684};
                15'd11179 : data_rom <= {16'd28771, 16'd15681};
                15'd11180 : data_rom <= {16'd28773, 16'd15678};
                15'd11181 : data_rom <= {16'd28774, 16'd15676};
                15'd11182 : data_rom <= {16'd28776, 16'd15673};
                15'd11183 : data_rom <= {16'd28777, 16'd15670};
                15'd11184 : data_rom <= {16'd28779, 16'd15667};
                15'd11185 : data_rom <= {16'd28780, 16'd15665};
                15'd11186 : data_rom <= {16'd28782, 16'd15662};
                15'd11187 : data_rom <= {16'd28783, 16'd15659};
                15'd11188 : data_rom <= {16'd28785, 16'd15656};
                15'd11189 : data_rom <= {16'd28786, 16'd15654};
                15'd11190 : data_rom <= {16'd28788, 16'd15651};
                15'd11191 : data_rom <= {16'd28789, 16'd15648};
                15'd11192 : data_rom <= {16'd28791, 16'd15645};
                15'd11193 : data_rom <= {16'd28792, 16'd15643};
                15'd11194 : data_rom <= {16'd28794, 16'd15640};
                15'd11195 : data_rom <= {16'd28795, 16'd15637};
                15'd11196 : data_rom <= {16'd28797, 16'd15634};
                15'd11197 : data_rom <= {16'd28798, 16'd15632};
                15'd11198 : data_rom <= {16'd28800, 16'd15629};
                15'd11199 : data_rom <= {16'd28801, 16'd15626};
                15'd11200 : data_rom <= {16'd28803, 16'd15623};
                15'd11201 : data_rom <= {16'd28804, 16'd15621};
                15'd11202 : data_rom <= {16'd28806, 16'd15618};
                15'd11203 : data_rom <= {16'd28807, 16'd15615};
                15'd11204 : data_rom <= {16'd28809, 16'd15612};
                15'd11205 : data_rom <= {16'd28810, 16'd15609};
                15'd11206 : data_rom <= {16'd28812, 16'd15607};
                15'd11207 : data_rom <= {16'd28813, 16'd15604};
                15'd11208 : data_rom <= {16'd28815, 16'd15601};
                15'd11209 : data_rom <= {16'd28816, 16'd15598};
                15'd11210 : data_rom <= {16'd28818, 16'd15596};
                15'd11211 : data_rom <= {16'd28819, 16'd15593};
                15'd11212 : data_rom <= {16'd28821, 16'd15590};
                15'd11213 : data_rom <= {16'd28822, 16'd15587};
                15'd11214 : data_rom <= {16'd28824, 16'd15585};
                15'd11215 : data_rom <= {16'd28825, 16'd15582};
                15'd11216 : data_rom <= {16'd28827, 16'd15579};
                15'd11217 : data_rom <= {16'd28828, 16'd15576};
                15'd11218 : data_rom <= {16'd28830, 16'd15574};
                15'd11219 : data_rom <= {16'd28831, 16'd15571};
                15'd11220 : data_rom <= {16'd28833, 16'd15568};
                15'd11221 : data_rom <= {16'd28834, 16'd15565};
                15'd11222 : data_rom <= {16'd28836, 16'd15562};
                15'd11223 : data_rom <= {16'd28837, 16'd15560};
                15'd11224 : data_rom <= {16'd28839, 16'd15557};
                15'd11225 : data_rom <= {16'd28840, 16'd15554};
                15'd11226 : data_rom <= {16'd28842, 16'd15551};
                15'd11227 : data_rom <= {16'd28843, 16'd15549};
                15'd11228 : data_rom <= {16'd28845, 16'd15546};
                15'd11229 : data_rom <= {16'd28846, 16'd15543};
                15'd11230 : data_rom <= {16'd28848, 16'd15540};
                15'd11231 : data_rom <= {16'd28849, 16'd15538};
                15'd11232 : data_rom <= {16'd28851, 16'd15535};
                15'd11233 : data_rom <= {16'd28852, 16'd15532};
                15'd11234 : data_rom <= {16'd28854, 16'd15529};
                15'd11235 : data_rom <= {16'd28855, 16'd15527};
                15'd11236 : data_rom <= {16'd28857, 16'd15524};
                15'd11237 : data_rom <= {16'd28858, 16'd15521};
                15'd11238 : data_rom <= {16'd28860, 16'd15518};
                15'd11239 : data_rom <= {16'd28861, 16'd15515};
                15'd11240 : data_rom <= {16'd28863, 16'd15513};
                15'd11241 : data_rom <= {16'd28864, 16'd15510};
                15'd11242 : data_rom <= {16'd28866, 16'd15507};
                15'd11243 : data_rom <= {16'd28867, 16'd15504};
                15'd11244 : data_rom <= {16'd28869, 16'd15502};
                15'd11245 : data_rom <= {16'd28870, 16'd15499};
                15'd11246 : data_rom <= {16'd28872, 16'd15496};
                15'd11247 : data_rom <= {16'd28873, 16'd15493};
                15'd11248 : data_rom <= {16'd28875, 16'd15491};
                15'd11249 : data_rom <= {16'd28876, 16'd15488};
                15'd11250 : data_rom <= {16'd28878, 16'd15485};
                15'd11251 : data_rom <= {16'd28879, 16'd15482};
                15'd11252 : data_rom <= {16'd28880, 16'd15479};
                15'd11253 : data_rom <= {16'd28882, 16'd15477};
                15'd11254 : data_rom <= {16'd28883, 16'd15474};
                15'd11255 : data_rom <= {16'd28885, 16'd15471};
                15'd11256 : data_rom <= {16'd28886, 16'd15468};
                15'd11257 : data_rom <= {16'd28888, 16'd15466};
                15'd11258 : data_rom <= {16'd28889, 16'd15463};
                15'd11259 : data_rom <= {16'd28891, 16'd15460};
                15'd11260 : data_rom <= {16'd28892, 16'd15457};
                15'd11261 : data_rom <= {16'd28894, 16'd15455};
                15'd11262 : data_rom <= {16'd28895, 16'd15452};
                15'd11263 : data_rom <= {16'd28897, 16'd15449};
                15'd11264 : data_rom <= {16'd28898, 16'd15446};
                15'd11265 : data_rom <= {16'd28900, 16'd15443};
                15'd11266 : data_rom <= {16'd28901, 16'd15441};
                15'd11267 : data_rom <= {16'd28903, 16'd15438};
                15'd11268 : data_rom <= {16'd28904, 16'd15435};
                15'd11269 : data_rom <= {16'd28906, 16'd15432};
                15'd11270 : data_rom <= {16'd28907, 16'd15430};
                15'd11271 : data_rom <= {16'd28909, 16'd15427};
                15'd11272 : data_rom <= {16'd28910, 16'd15424};
                15'd11273 : data_rom <= {16'd28912, 16'd15421};
                15'd11274 : data_rom <= {16'd28913, 16'd15419};
                15'd11275 : data_rom <= {16'd28915, 16'd15416};
                15'd11276 : data_rom <= {16'd28916, 16'd15413};
                15'd11277 : data_rom <= {16'd28918, 16'd15410};
                15'd11278 : data_rom <= {16'd28919, 16'd15407};
                15'd11279 : data_rom <= {16'd28920, 16'd15405};
                15'd11280 : data_rom <= {16'd28922, 16'd15402};
                15'd11281 : data_rom <= {16'd28923, 16'd15399};
                15'd11282 : data_rom <= {16'd28925, 16'd15396};
                15'd11283 : data_rom <= {16'd28926, 16'd15394};
                15'd11284 : data_rom <= {16'd28928, 16'd15391};
                15'd11285 : data_rom <= {16'd28929, 16'd15388};
                15'd11286 : data_rom <= {16'd28931, 16'd15385};
                15'd11287 : data_rom <= {16'd28932, 16'd15382};
                15'd11288 : data_rom <= {16'd28934, 16'd15380};
                15'd11289 : data_rom <= {16'd28935, 16'd15377};
                15'd11290 : data_rom <= {16'd28937, 16'd15374};
                15'd11291 : data_rom <= {16'd28938, 16'd15371};
                15'd11292 : data_rom <= {16'd28940, 16'd15369};
                15'd11293 : data_rom <= {16'd28941, 16'd15366};
                15'd11294 : data_rom <= {16'd28943, 16'd15363};
                15'd11295 : data_rom <= {16'd28944, 16'd15360};
                15'd11296 : data_rom <= {16'd28946, 16'd15358};
                15'd11297 : data_rom <= {16'd28947, 16'd15355};
                15'd11298 : data_rom <= {16'd28948, 16'd15352};
                15'd11299 : data_rom <= {16'd28950, 16'd15349};
                15'd11300 : data_rom <= {16'd28951, 16'd15346};
                15'd11301 : data_rom <= {16'd28953, 16'd15344};
                15'd11302 : data_rom <= {16'd28954, 16'd15341};
                15'd11303 : data_rom <= {16'd28956, 16'd15338};
                15'd11304 : data_rom <= {16'd28957, 16'd15335};
                15'd11305 : data_rom <= {16'd28959, 16'd15333};
                15'd11306 : data_rom <= {16'd28960, 16'd15330};
                15'd11307 : data_rom <= {16'd28962, 16'd15327};
                15'd11308 : data_rom <= {16'd28963, 16'd15324};
                15'd11309 : data_rom <= {16'd28965, 16'd15321};
                15'd11310 : data_rom <= {16'd28966, 16'd15319};
                15'd11311 : data_rom <= {16'd28968, 16'd15316};
                15'd11312 : data_rom <= {16'd28969, 16'd15313};
                15'd11313 : data_rom <= {16'd28971, 16'd15310};
                15'd11314 : data_rom <= {16'd28972, 16'd15308};
                15'd11315 : data_rom <= {16'd28973, 16'd15305};
                15'd11316 : data_rom <= {16'd28975, 16'd15302};
                15'd11317 : data_rom <= {16'd28976, 16'd15299};
                15'd11318 : data_rom <= {16'd28978, 16'd15296};
                15'd11319 : data_rom <= {16'd28979, 16'd15294};
                15'd11320 : data_rom <= {16'd28981, 16'd15291};
                15'd11321 : data_rom <= {16'd28982, 16'd15288};
                15'd11322 : data_rom <= {16'd28984, 16'd15285};
                15'd11323 : data_rom <= {16'd28985, 16'd15283};
                15'd11324 : data_rom <= {16'd28987, 16'd15280};
                15'd11325 : data_rom <= {16'd28988, 16'd15277};
                15'd11326 : data_rom <= {16'd28990, 16'd15274};
                15'd11327 : data_rom <= {16'd28991, 16'd15271};
                15'd11328 : data_rom <= {16'd28993, 16'd15269};
                15'd11329 : data_rom <= {16'd28994, 16'd15266};
                15'd11330 : data_rom <= {16'd28995, 16'd15263};
                15'd11331 : data_rom <= {16'd28997, 16'd15260};
                15'd11332 : data_rom <= {16'd28998, 16'd15258};
                15'd11333 : data_rom <= {16'd29000, 16'd15255};
                15'd11334 : data_rom <= {16'd29001, 16'd15252};
                15'd11335 : data_rom <= {16'd29003, 16'd15249};
                15'd11336 : data_rom <= {16'd29004, 16'd15246};
                15'd11337 : data_rom <= {16'd29006, 16'd15244};
                15'd11338 : data_rom <= {16'd29007, 16'd15241};
                15'd11339 : data_rom <= {16'd29009, 16'd15238};
                15'd11340 : data_rom <= {16'd29010, 16'd15235};
                15'd11341 : data_rom <= {16'd29012, 16'd15233};
                15'd11342 : data_rom <= {16'd29013, 16'd15230};
                15'd11343 : data_rom <= {16'd29014, 16'd15227};
                15'd11344 : data_rom <= {16'd29016, 16'd15224};
                15'd11345 : data_rom <= {16'd29017, 16'd15221};
                15'd11346 : data_rom <= {16'd29019, 16'd15219};
                15'd11347 : data_rom <= {16'd29020, 16'd15216};
                15'd11348 : data_rom <= {16'd29022, 16'd15213};
                15'd11349 : data_rom <= {16'd29023, 16'd15210};
                15'd11350 : data_rom <= {16'd29025, 16'd15207};
                15'd11351 : data_rom <= {16'd29026, 16'd15205};
                15'd11352 : data_rom <= {16'd29028, 16'd15202};
                15'd11353 : data_rom <= {16'd29029, 16'd15199};
                15'd11354 : data_rom <= {16'd29030, 16'd15196};
                15'd11355 : data_rom <= {16'd29032, 16'd15194};
                15'd11356 : data_rom <= {16'd29033, 16'd15191};
                15'd11357 : data_rom <= {16'd29035, 16'd15188};
                15'd11358 : data_rom <= {16'd29036, 16'd15185};
                15'd11359 : data_rom <= {16'd29038, 16'd15182};
                15'd11360 : data_rom <= {16'd29039, 16'd15180};
                15'd11361 : data_rom <= {16'd29041, 16'd15177};
                15'd11362 : data_rom <= {16'd29042, 16'd15174};
                15'd11363 : data_rom <= {16'd29044, 16'd15171};
                15'd11364 : data_rom <= {16'd29045, 16'd15168};
                15'd11365 : data_rom <= {16'd29046, 16'd15166};
                15'd11366 : data_rom <= {16'd29048, 16'd15163};
                15'd11367 : data_rom <= {16'd29049, 16'd15160};
                15'd11368 : data_rom <= {16'd29051, 16'd15157};
                15'd11369 : data_rom <= {16'd29052, 16'd15155};
                15'd11370 : data_rom <= {16'd29054, 16'd15152};
                15'd11371 : data_rom <= {16'd29055, 16'd15149};
                15'd11372 : data_rom <= {16'd29057, 16'd15146};
                15'd11373 : data_rom <= {16'd29058, 16'd15143};
                15'd11374 : data_rom <= {16'd29060, 16'd15141};
                15'd11375 : data_rom <= {16'd29061, 16'd15138};
                15'd11376 : data_rom <= {16'd29062, 16'd15135};
                15'd11377 : data_rom <= {16'd29064, 16'd15132};
                15'd11378 : data_rom <= {16'd29065, 16'd15129};
                15'd11379 : data_rom <= {16'd29067, 16'd15127};
                15'd11380 : data_rom <= {16'd29068, 16'd15124};
                15'd11381 : data_rom <= {16'd29070, 16'd15121};
                15'd11382 : data_rom <= {16'd29071, 16'd15118};
                15'd11383 : data_rom <= {16'd29073, 16'd15116};
                15'd11384 : data_rom <= {16'd29074, 16'd15113};
                15'd11385 : data_rom <= {16'd29076, 16'd15110};
                15'd11386 : data_rom <= {16'd29077, 16'd15107};
                15'd11387 : data_rom <= {16'd29078, 16'd15104};
                15'd11388 : data_rom <= {16'd29080, 16'd15102};
                15'd11389 : data_rom <= {16'd29081, 16'd15099};
                15'd11390 : data_rom <= {16'd29083, 16'd15096};
                15'd11391 : data_rom <= {16'd29084, 16'd15093};
                15'd11392 : data_rom <= {16'd29086, 16'd15090};
                15'd11393 : data_rom <= {16'd29087, 16'd15088};
                15'd11394 : data_rom <= {16'd29089, 16'd15085};
                15'd11395 : data_rom <= {16'd29090, 16'd15082};
                15'd11396 : data_rom <= {16'd29091, 16'd15079};
                15'd11397 : data_rom <= {16'd29093, 16'd15077};
                15'd11398 : data_rom <= {16'd29094, 16'd15074};
                15'd11399 : data_rom <= {16'd29096, 16'd15071};
                15'd11400 : data_rom <= {16'd29097, 16'd15068};
                15'd11401 : data_rom <= {16'd29099, 16'd15065};
                15'd11402 : data_rom <= {16'd29100, 16'd15063};
                15'd11403 : data_rom <= {16'd29102, 16'd15060};
                15'd11404 : data_rom <= {16'd29103, 16'd15057};
                15'd11405 : data_rom <= {16'd29104, 16'd15054};
                15'd11406 : data_rom <= {16'd29106, 16'd15051};
                15'd11407 : data_rom <= {16'd29107, 16'd15049};
                15'd11408 : data_rom <= {16'd29109, 16'd15046};
                15'd11409 : data_rom <= {16'd29110, 16'd15043};
                15'd11410 : data_rom <= {16'd29112, 16'd15040};
                15'd11411 : data_rom <= {16'd29113, 16'd15037};
                15'd11412 : data_rom <= {16'd29115, 16'd15035};
                15'd11413 : data_rom <= {16'd29116, 16'd15032};
                15'd11414 : data_rom <= {16'd29117, 16'd15029};
                15'd11415 : data_rom <= {16'd29119, 16'd15026};
                15'd11416 : data_rom <= {16'd29120, 16'd15023};
                15'd11417 : data_rom <= {16'd29122, 16'd15021};
                15'd11418 : data_rom <= {16'd29123, 16'd15018};
                15'd11419 : data_rom <= {16'd29125, 16'd15015};
                15'd11420 : data_rom <= {16'd29126, 16'd15012};
                15'd11421 : data_rom <= {16'd29128, 16'd15010};
                15'd11422 : data_rom <= {16'd29129, 16'd15007};
                15'd11423 : data_rom <= {16'd29130, 16'd15004};
                15'd11424 : data_rom <= {16'd29132, 16'd15001};
                15'd11425 : data_rom <= {16'd29133, 16'd14998};
                15'd11426 : data_rom <= {16'd29135, 16'd14996};
                15'd11427 : data_rom <= {16'd29136, 16'd14993};
                15'd11428 : data_rom <= {16'd29138, 16'd14990};
                15'd11429 : data_rom <= {16'd29139, 16'd14987};
                15'd11430 : data_rom <= {16'd29140, 16'd14984};
                15'd11431 : data_rom <= {16'd29142, 16'd14982};
                15'd11432 : data_rom <= {16'd29143, 16'd14979};
                15'd11433 : data_rom <= {16'd29145, 16'd14976};
                15'd11434 : data_rom <= {16'd29146, 16'd14973};
                15'd11435 : data_rom <= {16'd29148, 16'd14970};
                15'd11436 : data_rom <= {16'd29149, 16'd14968};
                15'd11437 : data_rom <= {16'd29150, 16'd14965};
                15'd11438 : data_rom <= {16'd29152, 16'd14962};
                15'd11439 : data_rom <= {16'd29153, 16'd14959};
                15'd11440 : data_rom <= {16'd29155, 16'd14956};
                15'd11441 : data_rom <= {16'd29156, 16'd14954};
                15'd11442 : data_rom <= {16'd29158, 16'd14951};
                15'd11443 : data_rom <= {16'd29159, 16'd14948};
                15'd11444 : data_rom <= {16'd29161, 16'd14945};
                15'd11445 : data_rom <= {16'd29162, 16'd14942};
                15'd11446 : data_rom <= {16'd29163, 16'd14940};
                15'd11447 : data_rom <= {16'd29165, 16'd14937};
                15'd11448 : data_rom <= {16'd29166, 16'd14934};
                15'd11449 : data_rom <= {16'd29168, 16'd14931};
                15'd11450 : data_rom <= {16'd29169, 16'd14928};
                15'd11451 : data_rom <= {16'd29171, 16'd14926};
                15'd11452 : data_rom <= {16'd29172, 16'd14923};
                15'd11453 : data_rom <= {16'd29173, 16'd14920};
                15'd11454 : data_rom <= {16'd29175, 16'd14917};
                15'd11455 : data_rom <= {16'd29176, 16'd14915};
                15'd11456 : data_rom <= {16'd29178, 16'd14912};
                15'd11457 : data_rom <= {16'd29179, 16'd14909};
                15'd11458 : data_rom <= {16'd29181, 16'd14906};
                15'd11459 : data_rom <= {16'd29182, 16'd14903};
                15'd11460 : data_rom <= {16'd29183, 16'd14901};
                15'd11461 : data_rom <= {16'd29185, 16'd14898};
                15'd11462 : data_rom <= {16'd29186, 16'd14895};
                15'd11463 : data_rom <= {16'd29188, 16'd14892};
                15'd11464 : data_rom <= {16'd29189, 16'd14889};
                15'd11465 : data_rom <= {16'd29191, 16'd14887};
                15'd11466 : data_rom <= {16'd29192, 16'd14884};
                15'd11467 : data_rom <= {16'd29193, 16'd14881};
                15'd11468 : data_rom <= {16'd29195, 16'd14878};
                15'd11469 : data_rom <= {16'd29196, 16'd14875};
                15'd11470 : data_rom <= {16'd29198, 16'd14873};
                15'd11471 : data_rom <= {16'd29199, 16'd14870};
                15'd11472 : data_rom <= {16'd29201, 16'd14867};
                15'd11473 : data_rom <= {16'd29202, 16'd14864};
                15'd11474 : data_rom <= {16'd29203, 16'd14861};
                15'd11475 : data_rom <= {16'd29205, 16'd14859};
                15'd11476 : data_rom <= {16'd29206, 16'd14856};
                15'd11477 : data_rom <= {16'd29208, 16'd14853};
                15'd11478 : data_rom <= {16'd29209, 16'd14850};
                15'd11479 : data_rom <= {16'd29211, 16'd14847};
                15'd11480 : data_rom <= {16'd29212, 16'd14845};
                15'd11481 : data_rom <= {16'd29213, 16'd14842};
                15'd11482 : data_rom <= {16'd29215, 16'd14839};
                15'd11483 : data_rom <= {16'd29216, 16'd14836};
                15'd11484 : data_rom <= {16'd29218, 16'd14833};
                15'd11485 : data_rom <= {16'd29219, 16'd14831};
                15'd11486 : data_rom <= {16'd29220, 16'd14828};
                15'd11487 : data_rom <= {16'd29222, 16'd14825};
                15'd11488 : data_rom <= {16'd29223, 16'd14822};
                15'd11489 : data_rom <= {16'd29225, 16'd14819};
                15'd11490 : data_rom <= {16'd29226, 16'd14817};
                15'd11491 : data_rom <= {16'd29228, 16'd14814};
                15'd11492 : data_rom <= {16'd29229, 16'd14811};
                15'd11493 : data_rom <= {16'd29230, 16'd14808};
                15'd11494 : data_rom <= {16'd29232, 16'd14805};
                15'd11495 : data_rom <= {16'd29233, 16'd14803};
                15'd11496 : data_rom <= {16'd29235, 16'd14800};
                15'd11497 : data_rom <= {16'd29236, 16'd14797};
                15'd11498 : data_rom <= {16'd29238, 16'd14794};
                15'd11499 : data_rom <= {16'd29239, 16'd14791};
                15'd11500 : data_rom <= {16'd29240, 16'd14788};
                15'd11501 : data_rom <= {16'd29242, 16'd14786};
                15'd11502 : data_rom <= {16'd29243, 16'd14783};
                15'd11503 : data_rom <= {16'd29245, 16'd14780};
                15'd11504 : data_rom <= {16'd29246, 16'd14777};
                15'd11505 : data_rom <= {16'd29247, 16'd14774};
                15'd11506 : data_rom <= {16'd29249, 16'd14772};
                15'd11507 : data_rom <= {16'd29250, 16'd14769};
                15'd11508 : data_rom <= {16'd29252, 16'd14766};
                15'd11509 : data_rom <= {16'd29253, 16'd14763};
                15'd11510 : data_rom <= {16'd29255, 16'd14760};
                15'd11511 : data_rom <= {16'd29256, 16'd14758};
                15'd11512 : data_rom <= {16'd29257, 16'd14755};
                15'd11513 : data_rom <= {16'd29259, 16'd14752};
                15'd11514 : data_rom <= {16'd29260, 16'd14749};
                15'd11515 : data_rom <= {16'd29262, 16'd14746};
                15'd11516 : data_rom <= {16'd29263, 16'd14744};
                15'd11517 : data_rom <= {16'd29264, 16'd14741};
                15'd11518 : data_rom <= {16'd29266, 16'd14738};
                15'd11519 : data_rom <= {16'd29267, 16'd14735};
                15'd11520 : data_rom <= {16'd29269, 16'd14732};
                15'd11521 : data_rom <= {16'd29270, 16'd14730};
                15'd11522 : data_rom <= {16'd29271, 16'd14727};
                15'd11523 : data_rom <= {16'd29273, 16'd14724};
                15'd11524 : data_rom <= {16'd29274, 16'd14721};
                15'd11525 : data_rom <= {16'd29276, 16'd14718};
                15'd11526 : data_rom <= {16'd29277, 16'd14716};
                15'd11527 : data_rom <= {16'd29279, 16'd14713};
                15'd11528 : data_rom <= {16'd29280, 16'd14710};
                15'd11529 : data_rom <= {16'd29281, 16'd14707};
                15'd11530 : data_rom <= {16'd29283, 16'd14704};
                15'd11531 : data_rom <= {16'd29284, 16'd14702};
                15'd11532 : data_rom <= {16'd29286, 16'd14699};
                15'd11533 : data_rom <= {16'd29287, 16'd14696};
                15'd11534 : data_rom <= {16'd29288, 16'd14693};
                15'd11535 : data_rom <= {16'd29290, 16'd14690};
                15'd11536 : data_rom <= {16'd29291, 16'd14687};
                15'd11537 : data_rom <= {16'd29293, 16'd14685};
                15'd11538 : data_rom <= {16'd29294, 16'd14682};
                15'd11539 : data_rom <= {16'd29295, 16'd14679};
                15'd11540 : data_rom <= {16'd29297, 16'd14676};
                15'd11541 : data_rom <= {16'd29298, 16'd14673};
                15'd11542 : data_rom <= {16'd29300, 16'd14671};
                15'd11543 : data_rom <= {16'd29301, 16'd14668};
                15'd11544 : data_rom <= {16'd29302, 16'd14665};
                15'd11545 : data_rom <= {16'd29304, 16'd14662};
                15'd11546 : data_rom <= {16'd29305, 16'd14659};
                15'd11547 : data_rom <= {16'd29307, 16'd14657};
                15'd11548 : data_rom <= {16'd29308, 16'd14654};
                15'd11549 : data_rom <= {16'd29310, 16'd14651};
                15'd11550 : data_rom <= {16'd29311, 16'd14648};
                15'd11551 : data_rom <= {16'd29312, 16'd14645};
                15'd11552 : data_rom <= {16'd29314, 16'd14643};
                15'd11553 : data_rom <= {16'd29315, 16'd14640};
                15'd11554 : data_rom <= {16'd29317, 16'd14637};
                15'd11555 : data_rom <= {16'd29318, 16'd14634};
                15'd11556 : data_rom <= {16'd29319, 16'd14631};
                15'd11557 : data_rom <= {16'd29321, 16'd14628};
                15'd11558 : data_rom <= {16'd29322, 16'd14626};
                15'd11559 : data_rom <= {16'd29324, 16'd14623};
                15'd11560 : data_rom <= {16'd29325, 16'd14620};
                15'd11561 : data_rom <= {16'd29326, 16'd14617};
                15'd11562 : data_rom <= {16'd29328, 16'd14614};
                15'd11563 : data_rom <= {16'd29329, 16'd14612};
                15'd11564 : data_rom <= {16'd29331, 16'd14609};
                15'd11565 : data_rom <= {16'd29332, 16'd14606};
                15'd11566 : data_rom <= {16'd29333, 16'd14603};
                15'd11567 : data_rom <= {16'd29335, 16'd14600};
                15'd11568 : data_rom <= {16'd29336, 16'd14598};
                15'd11569 : data_rom <= {16'd29338, 16'd14595};
                15'd11570 : data_rom <= {16'd29339, 16'd14592};
                15'd11571 : data_rom <= {16'd29340, 16'd14589};
                15'd11572 : data_rom <= {16'd29342, 16'd14586};
                15'd11573 : data_rom <= {16'd29343, 16'd14583};
                15'd11574 : data_rom <= {16'd29345, 16'd14581};
                15'd11575 : data_rom <= {16'd29346, 16'd14578};
                15'd11576 : data_rom <= {16'd29347, 16'd14575};
                15'd11577 : data_rom <= {16'd29349, 16'd14572};
                15'd11578 : data_rom <= {16'd29350, 16'd14569};
                15'd11579 : data_rom <= {16'd29352, 16'd14567};
                15'd11580 : data_rom <= {16'd29353, 16'd14564};
                15'd11581 : data_rom <= {16'd29354, 16'd14561};
                15'd11582 : data_rom <= {16'd29356, 16'd14558};
                15'd11583 : data_rom <= {16'd29357, 16'd14555};
                15'd11584 : data_rom <= {16'd29359, 16'd14553};
                15'd11585 : data_rom <= {16'd29360, 16'd14550};
                15'd11586 : data_rom <= {16'd29361, 16'd14547};
                15'd11587 : data_rom <= {16'd29363, 16'd14544};
                15'd11588 : data_rom <= {16'd29364, 16'd14541};
                15'd11589 : data_rom <= {16'd29365, 16'd14538};
                15'd11590 : data_rom <= {16'd29367, 16'd14536};
                15'd11591 : data_rom <= {16'd29368, 16'd14533};
                15'd11592 : data_rom <= {16'd29370, 16'd14530};
                15'd11593 : data_rom <= {16'd29371, 16'd14527};
                15'd11594 : data_rom <= {16'd29372, 16'd14524};
                15'd11595 : data_rom <= {16'd29374, 16'd14522};
                15'd11596 : data_rom <= {16'd29375, 16'd14519};
                15'd11597 : data_rom <= {16'd29377, 16'd14516};
                15'd11598 : data_rom <= {16'd29378, 16'd14513};
                15'd11599 : data_rom <= {16'd29379, 16'd14510};
                15'd11600 : data_rom <= {16'd29381, 16'd14507};
                15'd11601 : data_rom <= {16'd29382, 16'd14505};
                15'd11602 : data_rom <= {16'd29384, 16'd14502};
                15'd11603 : data_rom <= {16'd29385, 16'd14499};
                15'd11604 : data_rom <= {16'd29386, 16'd14496};
                15'd11605 : data_rom <= {16'd29388, 16'd14493};
                15'd11606 : data_rom <= {16'd29389, 16'd14491};
                15'd11607 : data_rom <= {16'd29391, 16'd14488};
                15'd11608 : data_rom <= {16'd29392, 16'd14485};
                15'd11609 : data_rom <= {16'd29393, 16'd14482};
                15'd11610 : data_rom <= {16'd29395, 16'd14479};
                15'd11611 : data_rom <= {16'd29396, 16'd14476};
                15'd11612 : data_rom <= {16'd29397, 16'd14474};
                15'd11613 : data_rom <= {16'd29399, 16'd14471};
                15'd11614 : data_rom <= {16'd29400, 16'd14468};
                15'd11615 : data_rom <= {16'd29402, 16'd14465};
                15'd11616 : data_rom <= {16'd29403, 16'd14462};
                15'd11617 : data_rom <= {16'd29404, 16'd14460};
                15'd11618 : data_rom <= {16'd29406, 16'd14457};
                15'd11619 : data_rom <= {16'd29407, 16'd14454};
                15'd11620 : data_rom <= {16'd29409, 16'd14451};
                15'd11621 : data_rom <= {16'd29410, 16'd14448};
                15'd11622 : data_rom <= {16'd29411, 16'd14445};
                15'd11623 : data_rom <= {16'd29413, 16'd14443};
                15'd11624 : data_rom <= {16'd29414, 16'd14440};
                15'd11625 : data_rom <= {16'd29415, 16'd14437};
                15'd11626 : data_rom <= {16'd29417, 16'd14434};
                15'd11627 : data_rom <= {16'd29418, 16'd14431};
                15'd11628 : data_rom <= {16'd29420, 16'd14429};
                15'd11629 : data_rom <= {16'd29421, 16'd14426};
                15'd11630 : data_rom <= {16'd29422, 16'd14423};
                15'd11631 : data_rom <= {16'd29424, 16'd14420};
                15'd11632 : data_rom <= {16'd29425, 16'd14417};
                15'd11633 : data_rom <= {16'd29427, 16'd14414};
                15'd11634 : data_rom <= {16'd29428, 16'd14412};
                15'd11635 : data_rom <= {16'd29429, 16'd14409};
                15'd11636 : data_rom <= {16'd29431, 16'd14406};
                15'd11637 : data_rom <= {16'd29432, 16'd14403};
                15'd11638 : data_rom <= {16'd29433, 16'd14400};
                15'd11639 : data_rom <= {16'd29435, 16'd14398};
                15'd11640 : data_rom <= {16'd29436, 16'd14395};
                15'd11641 : data_rom <= {16'd29438, 16'd14392};
                15'd11642 : data_rom <= {16'd29439, 16'd14389};
                15'd11643 : data_rom <= {16'd29440, 16'd14386};
                15'd11644 : data_rom <= {16'd29442, 16'd14383};
                15'd11645 : data_rom <= {16'd29443, 16'd14381};
                15'd11646 : data_rom <= {16'd29444, 16'd14378};
                15'd11647 : data_rom <= {16'd29446, 16'd14375};
                15'd11648 : data_rom <= {16'd29447, 16'd14372};
                15'd11649 : data_rom <= {16'd29449, 16'd14369};
                15'd11650 : data_rom <= {16'd29450, 16'd14366};
                15'd11651 : data_rom <= {16'd29451, 16'd14364};
                15'd11652 : data_rom <= {16'd29453, 16'd14361};
                15'd11653 : data_rom <= {16'd29454, 16'd14358};
                15'd11654 : data_rom <= {16'd29456, 16'd14355};
                15'd11655 : data_rom <= {16'd29457, 16'd14352};
                15'd11656 : data_rom <= {16'd29458, 16'd14350};
                15'd11657 : data_rom <= {16'd29460, 16'd14347};
                15'd11658 : data_rom <= {16'd29461, 16'd14344};
                15'd11659 : data_rom <= {16'd29462, 16'd14341};
                15'd11660 : data_rom <= {16'd29464, 16'd14338};
                15'd11661 : data_rom <= {16'd29465, 16'd14335};
                15'd11662 : data_rom <= {16'd29467, 16'd14333};
                15'd11663 : data_rom <= {16'd29468, 16'd14330};
                15'd11664 : data_rom <= {16'd29469, 16'd14327};
                15'd11665 : data_rom <= {16'd29471, 16'd14324};
                15'd11666 : data_rom <= {16'd29472, 16'd14321};
                15'd11667 : data_rom <= {16'd29473, 16'd14318};
                15'd11668 : data_rom <= {16'd29475, 16'd14316};
                15'd11669 : data_rom <= {16'd29476, 16'd14313};
                15'd11670 : data_rom <= {16'd29477, 16'd14310};
                15'd11671 : data_rom <= {16'd29479, 16'd14307};
                15'd11672 : data_rom <= {16'd29480, 16'd14304};
                15'd11673 : data_rom <= {16'd29482, 16'd14301};
                15'd11674 : data_rom <= {16'd29483, 16'd14299};
                15'd11675 : data_rom <= {16'd29484, 16'd14296};
                15'd11676 : data_rom <= {16'd29486, 16'd14293};
                15'd11677 : data_rom <= {16'd29487, 16'd14290};
                15'd11678 : data_rom <= {16'd29488, 16'd14287};
                15'd11679 : data_rom <= {16'd29490, 16'd14285};
                15'd11680 : data_rom <= {16'd29491, 16'd14282};
                15'd11681 : data_rom <= {16'd29493, 16'd14279};
                15'd11682 : data_rom <= {16'd29494, 16'd14276};
                15'd11683 : data_rom <= {16'd29495, 16'd14273};
                15'd11684 : data_rom <= {16'd29497, 16'd14270};
                15'd11685 : data_rom <= {16'd29498, 16'd14268};
                15'd11686 : data_rom <= {16'd29499, 16'd14265};
                15'd11687 : data_rom <= {16'd29501, 16'd14262};
                15'd11688 : data_rom <= {16'd29502, 16'd14259};
                15'd11689 : data_rom <= {16'd29504, 16'd14256};
                15'd11690 : data_rom <= {16'd29505, 16'd14253};
                15'd11691 : data_rom <= {16'd29506, 16'd14251};
                15'd11692 : data_rom <= {16'd29508, 16'd14248};
                15'd11693 : data_rom <= {16'd29509, 16'd14245};
                15'd11694 : data_rom <= {16'd29510, 16'd14242};
                15'd11695 : data_rom <= {16'd29512, 16'd14239};
                15'd11696 : data_rom <= {16'd29513, 16'd14236};
                15'd11697 : data_rom <= {16'd29514, 16'd14234};
                15'd11698 : data_rom <= {16'd29516, 16'd14231};
                15'd11699 : data_rom <= {16'd29517, 16'd14228};
                15'd11700 : data_rom <= {16'd29519, 16'd14225};
                15'd11701 : data_rom <= {16'd29520, 16'd14222};
                15'd11702 : data_rom <= {16'd29521, 16'd14219};
                15'd11703 : data_rom <= {16'd29523, 16'd14217};
                15'd11704 : data_rom <= {16'd29524, 16'd14214};
                15'd11705 : data_rom <= {16'd29525, 16'd14211};
                15'd11706 : data_rom <= {16'd29527, 16'd14208};
                15'd11707 : data_rom <= {16'd29528, 16'd14205};
                15'd11708 : data_rom <= {16'd29529, 16'd14202};
                15'd11709 : data_rom <= {16'd29531, 16'd14200};
                15'd11710 : data_rom <= {16'd29532, 16'd14197};
                15'd11711 : data_rom <= {16'd29534, 16'd14194};
                15'd11712 : data_rom <= {16'd29535, 16'd14191};
                15'd11713 : data_rom <= {16'd29536, 16'd14188};
                15'd11714 : data_rom <= {16'd29538, 16'd14185};
                15'd11715 : data_rom <= {16'd29539, 16'd14183};
                15'd11716 : data_rom <= {16'd29540, 16'd14180};
                15'd11717 : data_rom <= {16'd29542, 16'd14177};
                15'd11718 : data_rom <= {16'd29543, 16'd14174};
                15'd11719 : data_rom <= {16'd29544, 16'd14171};
                15'd11720 : data_rom <= {16'd29546, 16'd14168};
                15'd11721 : data_rom <= {16'd29547, 16'd14166};
                15'd11722 : data_rom <= {16'd29548, 16'd14163};
                15'd11723 : data_rom <= {16'd29550, 16'd14160};
                15'd11724 : data_rom <= {16'd29551, 16'd14157};
                15'd11725 : data_rom <= {16'd29553, 16'd14154};
                15'd11726 : data_rom <= {16'd29554, 16'd14151};
                15'd11727 : data_rom <= {16'd29555, 16'd14149};
                15'd11728 : data_rom <= {16'd29557, 16'd14146};
                15'd11729 : data_rom <= {16'd29558, 16'd14143};
                15'd11730 : data_rom <= {16'd29559, 16'd14140};
                15'd11731 : data_rom <= {16'd29561, 16'd14137};
                15'd11732 : data_rom <= {16'd29562, 16'd14134};
                15'd11733 : data_rom <= {16'd29563, 16'd14132};
                15'd11734 : data_rom <= {16'd29565, 16'd14129};
                15'd11735 : data_rom <= {16'd29566, 16'd14126};
                15'd11736 : data_rom <= {16'd29567, 16'd14123};
                15'd11737 : data_rom <= {16'd29569, 16'd14120};
                15'd11738 : data_rom <= {16'd29570, 16'd14117};
                15'd11739 : data_rom <= {16'd29572, 16'd14115};
                15'd11740 : data_rom <= {16'd29573, 16'd14112};
                15'd11741 : data_rom <= {16'd29574, 16'd14109};
                15'd11742 : data_rom <= {16'd29576, 16'd14106};
                15'd11743 : data_rom <= {16'd29577, 16'd14103};
                15'd11744 : data_rom <= {16'd29578, 16'd14100};
                15'd11745 : data_rom <= {16'd29580, 16'd14098};
                15'd11746 : data_rom <= {16'd29581, 16'd14095};
                15'd11747 : data_rom <= {16'd29582, 16'd14092};
                15'd11748 : data_rom <= {16'd29584, 16'd14089};
                15'd11749 : data_rom <= {16'd29585, 16'd14086};
                15'd11750 : data_rom <= {16'd29586, 16'd14083};
                15'd11751 : data_rom <= {16'd29588, 16'd14081};
                15'd11752 : data_rom <= {16'd29589, 16'd14078};
                15'd11753 : data_rom <= {16'd29590, 16'd14075};
                15'd11754 : data_rom <= {16'd29592, 16'd14072};
                15'd11755 : data_rom <= {16'd29593, 16'd14069};
                15'd11756 : data_rom <= {16'd29594, 16'd14066};
                15'd11757 : data_rom <= {16'd29596, 16'd14064};
                15'd11758 : data_rom <= {16'd29597, 16'd14061};
                15'd11759 : data_rom <= {16'd29599, 16'd14058};
                15'd11760 : data_rom <= {16'd29600, 16'd14055};
                15'd11761 : data_rom <= {16'd29601, 16'd14052};
                15'd11762 : data_rom <= {16'd29603, 16'd14049};
                15'd11763 : data_rom <= {16'd29604, 16'd14047};
                15'd11764 : data_rom <= {16'd29605, 16'd14044};
                15'd11765 : data_rom <= {16'd29607, 16'd14041};
                15'd11766 : data_rom <= {16'd29608, 16'd14038};
                15'd11767 : data_rom <= {16'd29609, 16'd14035};
                15'd11768 : data_rom <= {16'd29611, 16'd14032};
                15'd11769 : data_rom <= {16'd29612, 16'd14030};
                15'd11770 : data_rom <= {16'd29613, 16'd14027};
                15'd11771 : data_rom <= {16'd29615, 16'd14024};
                15'd11772 : data_rom <= {16'd29616, 16'd14021};
                15'd11773 : data_rom <= {16'd29617, 16'd14018};
                15'd11774 : data_rom <= {16'd29619, 16'd14015};
                15'd11775 : data_rom <= {16'd29620, 16'd14012};
                15'd11776 : data_rom <= {16'd29621, 16'd14010};
                15'd11777 : data_rom <= {16'd29623, 16'd14007};
                15'd11778 : data_rom <= {16'd29624, 16'd14004};
                15'd11779 : data_rom <= {16'd29625, 16'd14001};
                15'd11780 : data_rom <= {16'd29627, 16'd13998};
                15'd11781 : data_rom <= {16'd29628, 16'd13995};
                15'd11782 : data_rom <= {16'd29629, 16'd13993};
                15'd11783 : data_rom <= {16'd29631, 16'd13990};
                15'd11784 : data_rom <= {16'd29632, 16'd13987};
                15'd11785 : data_rom <= {16'd29633, 16'd13984};
                15'd11786 : data_rom <= {16'd29635, 16'd13981};
                15'd11787 : data_rom <= {16'd29636, 16'd13978};
                15'd11788 : data_rom <= {16'd29638, 16'd13976};
                15'd11789 : data_rom <= {16'd29639, 16'd13973};
                15'd11790 : data_rom <= {16'd29640, 16'd13970};
                15'd11791 : data_rom <= {16'd29642, 16'd13967};
                15'd11792 : data_rom <= {16'd29643, 16'd13964};
                15'd11793 : data_rom <= {16'd29644, 16'd13961};
                15'd11794 : data_rom <= {16'd29646, 16'd13959};
                15'd11795 : data_rom <= {16'd29647, 16'd13956};
                15'd11796 : data_rom <= {16'd29648, 16'd13953};
                15'd11797 : data_rom <= {16'd29650, 16'd13950};
                15'd11798 : data_rom <= {16'd29651, 16'd13947};
                15'd11799 : data_rom <= {16'd29652, 16'd13944};
                15'd11800 : data_rom <= {16'd29654, 16'd13941};
                15'd11801 : data_rom <= {16'd29655, 16'd13939};
                15'd11802 : data_rom <= {16'd29656, 16'd13936};
                15'd11803 : data_rom <= {16'd29658, 16'd13933};
                15'd11804 : data_rom <= {16'd29659, 16'd13930};
                15'd11805 : data_rom <= {16'd29660, 16'd13927};
                15'd11806 : data_rom <= {16'd29662, 16'd13924};
                15'd11807 : data_rom <= {16'd29663, 16'd13922};
                15'd11808 : data_rom <= {16'd29664, 16'd13919};
                15'd11809 : data_rom <= {16'd29666, 16'd13916};
                15'd11810 : data_rom <= {16'd29667, 16'd13913};
                15'd11811 : data_rom <= {16'd29668, 16'd13910};
                15'd11812 : data_rom <= {16'd29670, 16'd13907};
                15'd11813 : data_rom <= {16'd29671, 16'd13904};
                15'd11814 : data_rom <= {16'd29672, 16'd13902};
                15'd11815 : data_rom <= {16'd29674, 16'd13899};
                15'd11816 : data_rom <= {16'd29675, 16'd13896};
                15'd11817 : data_rom <= {16'd29676, 16'd13893};
                15'd11818 : data_rom <= {16'd29678, 16'd13890};
                15'd11819 : data_rom <= {16'd29679, 16'd13887};
                15'd11820 : data_rom <= {16'd29680, 16'd13885};
                15'd11821 : data_rom <= {16'd29682, 16'd13882};
                15'd11822 : data_rom <= {16'd29683, 16'd13879};
                15'd11823 : data_rom <= {16'd29684, 16'd13876};
                15'd11824 : data_rom <= {16'd29686, 16'd13873};
                15'd11825 : data_rom <= {16'd29687, 16'd13870};
                15'd11826 : data_rom <= {16'd29688, 16'd13867};
                15'd11827 : data_rom <= {16'd29690, 16'd13865};
                15'd11828 : data_rom <= {16'd29691, 16'd13862};
                15'd11829 : data_rom <= {16'd29692, 16'd13859};
                15'd11830 : data_rom <= {16'd29694, 16'd13856};
                15'd11831 : data_rom <= {16'd29695, 16'd13853};
                15'd11832 : data_rom <= {16'd29696, 16'd13850};
                15'd11833 : data_rom <= {16'd29698, 16'd13848};
                15'd11834 : data_rom <= {16'd29699, 16'd13845};
                15'd11835 : data_rom <= {16'd29700, 16'd13842};
                15'd11836 : data_rom <= {16'd29702, 16'd13839};
                15'd11837 : data_rom <= {16'd29703, 16'd13836};
                15'd11838 : data_rom <= {16'd29704, 16'd13833};
                15'd11839 : data_rom <= {16'd29705, 16'd13830};
                15'd11840 : data_rom <= {16'd29707, 16'd13828};
                15'd11841 : data_rom <= {16'd29708, 16'd13825};
                15'd11842 : data_rom <= {16'd29709, 16'd13822};
                15'd11843 : data_rom <= {16'd29711, 16'd13819};
                15'd11844 : data_rom <= {16'd29712, 16'd13816};
                15'd11845 : data_rom <= {16'd29713, 16'd13813};
                15'd11846 : data_rom <= {16'd29715, 16'd13811};
                15'd11847 : data_rom <= {16'd29716, 16'd13808};
                15'd11848 : data_rom <= {16'd29717, 16'd13805};
                15'd11849 : data_rom <= {16'd29719, 16'd13802};
                15'd11850 : data_rom <= {16'd29720, 16'd13799};
                15'd11851 : data_rom <= {16'd29721, 16'd13796};
                15'd11852 : data_rom <= {16'd29723, 16'd13793};
                15'd11853 : data_rom <= {16'd29724, 16'd13791};
                15'd11854 : data_rom <= {16'd29725, 16'd13788};
                15'd11855 : data_rom <= {16'd29727, 16'd13785};
                15'd11856 : data_rom <= {16'd29728, 16'd13782};
                15'd11857 : data_rom <= {16'd29729, 16'd13779};
                15'd11858 : data_rom <= {16'd29731, 16'd13776};
                15'd11859 : data_rom <= {16'd29732, 16'd13773};
                15'd11860 : data_rom <= {16'd29733, 16'd13771};
                15'd11861 : data_rom <= {16'd29735, 16'd13768};
                15'd11862 : data_rom <= {16'd29736, 16'd13765};
                15'd11863 : data_rom <= {16'd29737, 16'd13762};
                15'd11864 : data_rom <= {16'd29739, 16'd13759};
                15'd11865 : data_rom <= {16'd29740, 16'd13756};
                15'd11866 : data_rom <= {16'd29741, 16'd13754};
                15'd11867 : data_rom <= {16'd29743, 16'd13751};
                15'd11868 : data_rom <= {16'd29744, 16'd13748};
                15'd11869 : data_rom <= {16'd29745, 16'd13745};
                15'd11870 : data_rom <= {16'd29746, 16'd13742};
                15'd11871 : data_rom <= {16'd29748, 16'd13739};
                15'd11872 : data_rom <= {16'd29749, 16'd13736};
                15'd11873 : data_rom <= {16'd29750, 16'd13734};
                15'd11874 : data_rom <= {16'd29752, 16'd13731};
                15'd11875 : data_rom <= {16'd29753, 16'd13728};
                15'd11876 : data_rom <= {16'd29754, 16'd13725};
                15'd11877 : data_rom <= {16'd29756, 16'd13722};
                15'd11878 : data_rom <= {16'd29757, 16'd13719};
                15'd11879 : data_rom <= {16'd29758, 16'd13716};
                15'd11880 : data_rom <= {16'd29760, 16'd13714};
                15'd11881 : data_rom <= {16'd29761, 16'd13711};
                15'd11882 : data_rom <= {16'd29762, 16'd13708};
                15'd11883 : data_rom <= {16'd29764, 16'd13705};
                15'd11884 : data_rom <= {16'd29765, 16'd13702};
                15'd11885 : data_rom <= {16'd29766, 16'd13699};
                15'd11886 : data_rom <= {16'd29768, 16'd13696};
                15'd11887 : data_rom <= {16'd29769, 16'd13694};
                15'd11888 : data_rom <= {16'd29770, 16'd13691};
                15'd11889 : data_rom <= {16'd29771, 16'd13688};
                15'd11890 : data_rom <= {16'd29773, 16'd13685};
                15'd11891 : data_rom <= {16'd29774, 16'd13682};
                15'd11892 : data_rom <= {16'd29775, 16'd13679};
                15'd11893 : data_rom <= {16'd29777, 16'd13677};
                15'd11894 : data_rom <= {16'd29778, 16'd13674};
                15'd11895 : data_rom <= {16'd29779, 16'd13671};
                15'd11896 : data_rom <= {16'd29781, 16'd13668};
                15'd11897 : data_rom <= {16'd29782, 16'd13665};
                15'd11898 : data_rom <= {16'd29783, 16'd13662};
                15'd11899 : data_rom <= {16'd29785, 16'd13659};
                15'd11900 : data_rom <= {16'd29786, 16'd13657};
                15'd11901 : data_rom <= {16'd29787, 16'd13654};
                15'd11902 : data_rom <= {16'd29788, 16'd13651};
                15'd11903 : data_rom <= {16'd29790, 16'd13648};
                15'd11904 : data_rom <= {16'd29791, 16'd13645};
                15'd11905 : data_rom <= {16'd29792, 16'd13642};
                15'd11906 : data_rom <= {16'd29794, 16'd13639};
                15'd11907 : data_rom <= {16'd29795, 16'd13637};
                15'd11908 : data_rom <= {16'd29796, 16'd13634};
                15'd11909 : data_rom <= {16'd29798, 16'd13631};
                15'd11910 : data_rom <= {16'd29799, 16'd13628};
                15'd11911 : data_rom <= {16'd29800, 16'd13625};
                15'd11912 : data_rom <= {16'd29802, 16'd13622};
                15'd11913 : data_rom <= {16'd29803, 16'd13619};
                15'd11914 : data_rom <= {16'd29804, 16'd13617};
                15'd11915 : data_rom <= {16'd29805, 16'd13614};
                15'd11916 : data_rom <= {16'd29807, 16'd13611};
                15'd11917 : data_rom <= {16'd29808, 16'd13608};
                15'd11918 : data_rom <= {16'd29809, 16'd13605};
                15'd11919 : data_rom <= {16'd29811, 16'd13602};
                15'd11920 : data_rom <= {16'd29812, 16'd13599};
                15'd11921 : data_rom <= {16'd29813, 16'd13597};
                15'd11922 : data_rom <= {16'd29815, 16'd13594};
                15'd11923 : data_rom <= {16'd29816, 16'd13591};
                15'd11924 : data_rom <= {16'd29817, 16'd13588};
                15'd11925 : data_rom <= {16'd29819, 16'd13585};
                15'd11926 : data_rom <= {16'd29820, 16'd13582};
                15'd11927 : data_rom <= {16'd29821, 16'd13579};
                15'd11928 : data_rom <= {16'd29822, 16'd13577};
                15'd11929 : data_rom <= {16'd29824, 16'd13574};
                15'd11930 : data_rom <= {16'd29825, 16'd13571};
                15'd11931 : data_rom <= {16'd29826, 16'd13568};
                15'd11932 : data_rom <= {16'd29828, 16'd13565};
                15'd11933 : data_rom <= {16'd29829, 16'd13562};
                15'd11934 : data_rom <= {16'd29830, 16'd13559};
                15'd11935 : data_rom <= {16'd29832, 16'd13556};
                15'd11936 : data_rom <= {16'd29833, 16'd13554};
                15'd11937 : data_rom <= {16'd29834, 16'd13551};
                15'd11938 : data_rom <= {16'd29835, 16'd13548};
                15'd11939 : data_rom <= {16'd29837, 16'd13545};
                15'd11940 : data_rom <= {16'd29838, 16'd13542};
                15'd11941 : data_rom <= {16'd29839, 16'd13539};
                15'd11942 : data_rom <= {16'd29841, 16'd13536};
                15'd11943 : data_rom <= {16'd29842, 16'd13534};
                15'd11944 : data_rom <= {16'd29843, 16'd13531};
                15'd11945 : data_rom <= {16'd29845, 16'd13528};
                15'd11946 : data_rom <= {16'd29846, 16'd13525};
                15'd11947 : data_rom <= {16'd29847, 16'd13522};
                15'd11948 : data_rom <= {16'd29848, 16'd13519};
                15'd11949 : data_rom <= {16'd29850, 16'd13516};
                15'd11950 : data_rom <= {16'd29851, 16'd13514};
                15'd11951 : data_rom <= {16'd29852, 16'd13511};
                15'd11952 : data_rom <= {16'd29854, 16'd13508};
                15'd11953 : data_rom <= {16'd29855, 16'd13505};
                15'd11954 : data_rom <= {16'd29856, 16'd13502};
                15'd11955 : data_rom <= {16'd29857, 16'd13499};
                15'd11956 : data_rom <= {16'd29859, 16'd13496};
                15'd11957 : data_rom <= {16'd29860, 16'd13494};
                15'd11958 : data_rom <= {16'd29861, 16'd13491};
                15'd11959 : data_rom <= {16'd29863, 16'd13488};
                15'd11960 : data_rom <= {16'd29864, 16'd13485};
                15'd11961 : data_rom <= {16'd29865, 16'd13482};
                15'd11962 : data_rom <= {16'd29867, 16'd13479};
                15'd11963 : data_rom <= {16'd29868, 16'd13476};
                15'd11964 : data_rom <= {16'd29869, 16'd13473};
                15'd11965 : data_rom <= {16'd29870, 16'd13471};
                15'd11966 : data_rom <= {16'd29872, 16'd13468};
                15'd11967 : data_rom <= {16'd29873, 16'd13465};
                15'd11968 : data_rom <= {16'd29874, 16'd13462};
                15'd11969 : data_rom <= {16'd29876, 16'd13459};
                15'd11970 : data_rom <= {16'd29877, 16'd13456};
                15'd11971 : data_rom <= {16'd29878, 16'd13453};
                15'd11972 : data_rom <= {16'd29879, 16'd13451};
                15'd11973 : data_rom <= {16'd29881, 16'd13448};
                15'd11974 : data_rom <= {16'd29882, 16'd13445};
                15'd11975 : data_rom <= {16'd29883, 16'd13442};
                15'd11976 : data_rom <= {16'd29885, 16'd13439};
                15'd11977 : data_rom <= {16'd29886, 16'd13436};
                15'd11978 : data_rom <= {16'd29887, 16'd13433};
                15'd11979 : data_rom <= {16'd29888, 16'd13431};
                15'd11980 : data_rom <= {16'd29890, 16'd13428};
                15'd11981 : data_rom <= {16'd29891, 16'd13425};
                15'd11982 : data_rom <= {16'd29892, 16'd13422};
                15'd11983 : data_rom <= {16'd29894, 16'd13419};
                15'd11984 : data_rom <= {16'd29895, 16'd13416};
                15'd11985 : data_rom <= {16'd29896, 16'd13413};
                15'd11986 : data_rom <= {16'd29897, 16'd13410};
                15'd11987 : data_rom <= {16'd29899, 16'd13408};
                15'd11988 : data_rom <= {16'd29900, 16'd13405};
                15'd11989 : data_rom <= {16'd29901, 16'd13402};
                15'd11990 : data_rom <= {16'd29903, 16'd13399};
                15'd11991 : data_rom <= {16'd29904, 16'd13396};
                15'd11992 : data_rom <= {16'd29905, 16'd13393};
                15'd11993 : data_rom <= {16'd29906, 16'd13390};
                15'd11994 : data_rom <= {16'd29908, 16'd13388};
                15'd11995 : data_rom <= {16'd29909, 16'd13385};
                15'd11996 : data_rom <= {16'd29910, 16'd13382};
                15'd11997 : data_rom <= {16'd29912, 16'd13379};
                15'd11998 : data_rom <= {16'd29913, 16'd13376};
                15'd11999 : data_rom <= {16'd29914, 16'd13373};
                15'd12000 : data_rom <= {16'd29915, 16'd13370};
                15'd12001 : data_rom <= {16'd29917, 16'd13367};
                15'd12002 : data_rom <= {16'd29918, 16'd13365};
                15'd12003 : data_rom <= {16'd29919, 16'd13362};
                15'd12004 : data_rom <= {16'd29921, 16'd13359};
                15'd12005 : data_rom <= {16'd29922, 16'd13356};
                15'd12006 : data_rom <= {16'd29923, 16'd13353};
                15'd12007 : data_rom <= {16'd29924, 16'd13350};
                15'd12008 : data_rom <= {16'd29926, 16'd13347};
                15'd12009 : data_rom <= {16'd29927, 16'd13345};
                15'd12010 : data_rom <= {16'd29928, 16'd13342};
                15'd12011 : data_rom <= {16'd29930, 16'd13339};
                15'd12012 : data_rom <= {16'd29931, 16'd13336};
                15'd12013 : data_rom <= {16'd29932, 16'd13333};
                15'd12014 : data_rom <= {16'd29933, 16'd13330};
                15'd12015 : data_rom <= {16'd29935, 16'd13327};
                15'd12016 : data_rom <= {16'd29936, 16'd13324};
                15'd12017 : data_rom <= {16'd29937, 16'd13322};
                15'd12018 : data_rom <= {16'd29938, 16'd13319};
                15'd12019 : data_rom <= {16'd29940, 16'd13316};
                15'd12020 : data_rom <= {16'd29941, 16'd13313};
                15'd12021 : data_rom <= {16'd29942, 16'd13310};
                15'd12022 : data_rom <= {16'd29944, 16'd13307};
                15'd12023 : data_rom <= {16'd29945, 16'd13304};
                15'd12024 : data_rom <= {16'd29946, 16'd13301};
                15'd12025 : data_rom <= {16'd29947, 16'd13299};
                15'd12026 : data_rom <= {16'd29949, 16'd13296};
                15'd12027 : data_rom <= {16'd29950, 16'd13293};
                15'd12028 : data_rom <= {16'd29951, 16'd13290};
                15'd12029 : data_rom <= {16'd29952, 16'd13287};
                15'd12030 : data_rom <= {16'd29954, 16'd13284};
                15'd12031 : data_rom <= {16'd29955, 16'd13281};
                15'd12032 : data_rom <= {16'd29956, 16'd13278};
                15'd12033 : data_rom <= {16'd29958, 16'd13276};
                15'd12034 : data_rom <= {16'd29959, 16'd13273};
                15'd12035 : data_rom <= {16'd29960, 16'd13270};
                15'd12036 : data_rom <= {16'd29961, 16'd13267};
                15'd12037 : data_rom <= {16'd29963, 16'd13264};
                15'd12038 : data_rom <= {16'd29964, 16'd13261};
                15'd12039 : data_rom <= {16'd29965, 16'd13258};
                15'd12040 : data_rom <= {16'd29966, 16'd13255};
                15'd12041 : data_rom <= {16'd29968, 16'd13253};
                15'd12042 : data_rom <= {16'd29969, 16'd13250};
                15'd12043 : data_rom <= {16'd29970, 16'd13247};
                15'd12044 : data_rom <= {16'd29972, 16'd13244};
                15'd12045 : data_rom <= {16'd29973, 16'd13241};
                15'd12046 : data_rom <= {16'd29974, 16'd13238};
                15'd12047 : data_rom <= {16'd29975, 16'd13235};
                15'd12048 : data_rom <= {16'd29977, 16'd13233};
                15'd12049 : data_rom <= {16'd29978, 16'd13230};
                15'd12050 : data_rom <= {16'd29979, 16'd13227};
                15'd12051 : data_rom <= {16'd29980, 16'd13224};
                15'd12052 : data_rom <= {16'd29982, 16'd13221};
                15'd12053 : data_rom <= {16'd29983, 16'd13218};
                15'd12054 : data_rom <= {16'd29984, 16'd13215};
                15'd12055 : data_rom <= {16'd29986, 16'd13212};
                15'd12056 : data_rom <= {16'd29987, 16'd13210};
                15'd12057 : data_rom <= {16'd29988, 16'd13207};
                15'd12058 : data_rom <= {16'd29989, 16'd13204};
                15'd12059 : data_rom <= {16'd29991, 16'd13201};
                15'd12060 : data_rom <= {16'd29992, 16'd13198};
                15'd12061 : data_rom <= {16'd29993, 16'd13195};
                15'd12062 : data_rom <= {16'd29994, 16'd13192};
                15'd12063 : data_rom <= {16'd29996, 16'd13189};
                15'd12064 : data_rom <= {16'd29997, 16'd13187};
                15'd12065 : data_rom <= {16'd29998, 16'd13184};
                15'd12066 : data_rom <= {16'd29999, 16'd13181};
                15'd12067 : data_rom <= {16'd30001, 16'd13178};
                15'd12068 : data_rom <= {16'd30002, 16'd13175};
                15'd12069 : data_rom <= {16'd30003, 16'd13172};
                15'd12070 : data_rom <= {16'd30004, 16'd13169};
                15'd12071 : data_rom <= {16'd30006, 16'd13166};
                15'd12072 : data_rom <= {16'd30007, 16'd13163};
                15'd12073 : data_rom <= {16'd30008, 16'd13161};
                15'd12074 : data_rom <= {16'd30010, 16'd13158};
                15'd12075 : data_rom <= {16'd30011, 16'd13155};
                15'd12076 : data_rom <= {16'd30012, 16'd13152};
                15'd12077 : data_rom <= {16'd30013, 16'd13149};
                15'd12078 : data_rom <= {16'd30015, 16'd13146};
                15'd12079 : data_rom <= {16'd30016, 16'd13143};
                15'd12080 : data_rom <= {16'd30017, 16'd13140};
                15'd12081 : data_rom <= {16'd30018, 16'd13138};
                15'd12082 : data_rom <= {16'd30020, 16'd13135};
                15'd12083 : data_rom <= {16'd30021, 16'd13132};
                15'd12084 : data_rom <= {16'd30022, 16'd13129};
                15'd12085 : data_rom <= {16'd30023, 16'd13126};
                15'd12086 : data_rom <= {16'd30025, 16'd13123};
                15'd12087 : data_rom <= {16'd30026, 16'd13120};
                15'd12088 : data_rom <= {16'd30027, 16'd13117};
                15'd12089 : data_rom <= {16'd30028, 16'd13115};
                15'd12090 : data_rom <= {16'd30030, 16'd13112};
                15'd12091 : data_rom <= {16'd30031, 16'd13109};
                15'd12092 : data_rom <= {16'd30032, 16'd13106};
                15'd12093 : data_rom <= {16'd30033, 16'd13103};
                15'd12094 : data_rom <= {16'd30035, 16'd13100};
                15'd12095 : data_rom <= {16'd30036, 16'd13097};
                15'd12096 : data_rom <= {16'd30037, 16'd13094};
                15'd12097 : data_rom <= {16'd30038, 16'd13092};
                15'd12098 : data_rom <= {16'd30040, 16'd13089};
                15'd12099 : data_rom <= {16'd30041, 16'd13086};
                15'd12100 : data_rom <= {16'd30042, 16'd13083};
                15'd12101 : data_rom <= {16'd30043, 16'd13080};
                15'd12102 : data_rom <= {16'd30045, 16'd13077};
                15'd12103 : data_rom <= {16'd30046, 16'd13074};
                15'd12104 : data_rom <= {16'd30047, 16'd13071};
                15'd12105 : data_rom <= {16'd30049, 16'd13068};
                15'd12106 : data_rom <= {16'd30050, 16'd13066};
                15'd12107 : data_rom <= {16'd30051, 16'd13063};
                15'd12108 : data_rom <= {16'd30052, 16'd13060};
                15'd12109 : data_rom <= {16'd30054, 16'd13057};
                15'd12110 : data_rom <= {16'd30055, 16'd13054};
                15'd12111 : data_rom <= {16'd30056, 16'd13051};
                15'd12112 : data_rom <= {16'd30057, 16'd13048};
                15'd12113 : data_rom <= {16'd30059, 16'd13045};
                15'd12114 : data_rom <= {16'd30060, 16'd13043};
                15'd12115 : data_rom <= {16'd30061, 16'd13040};
                15'd12116 : data_rom <= {16'd30062, 16'd13037};
                15'd12117 : data_rom <= {16'd30064, 16'd13034};
                15'd12118 : data_rom <= {16'd30065, 16'd13031};
                15'd12119 : data_rom <= {16'd30066, 16'd13028};
                15'd12120 : data_rom <= {16'd30067, 16'd13025};
                15'd12121 : data_rom <= {16'd30069, 16'd13022};
                15'd12122 : data_rom <= {16'd30070, 16'd13020};
                15'd12123 : data_rom <= {16'd30071, 16'd13017};
                15'd12124 : data_rom <= {16'd30072, 16'd13014};
                15'd12125 : data_rom <= {16'd30074, 16'd13011};
                15'd12126 : data_rom <= {16'd30075, 16'd13008};
                15'd12127 : data_rom <= {16'd30076, 16'd13005};
                15'd12128 : data_rom <= {16'd30077, 16'd13002};
                15'd12129 : data_rom <= {16'd30079, 16'd12999};
                15'd12130 : data_rom <= {16'd30080, 16'd12996};
                15'd12131 : data_rom <= {16'd30081, 16'd12994};
                15'd12132 : data_rom <= {16'd30082, 16'd12991};
                15'd12133 : data_rom <= {16'd30083, 16'd12988};
                15'd12134 : data_rom <= {16'd30085, 16'd12985};
                15'd12135 : data_rom <= {16'd30086, 16'd12982};
                15'd12136 : data_rom <= {16'd30087, 16'd12979};
                15'd12137 : data_rom <= {16'd30088, 16'd12976};
                15'd12138 : data_rom <= {16'd30090, 16'd12973};
                15'd12139 : data_rom <= {16'd30091, 16'd12970};
                15'd12140 : data_rom <= {16'd30092, 16'd12968};
                15'd12141 : data_rom <= {16'd30093, 16'd12965};
                15'd12142 : data_rom <= {16'd30095, 16'd12962};
                15'd12143 : data_rom <= {16'd30096, 16'd12959};
                15'd12144 : data_rom <= {16'd30097, 16'd12956};
                15'd12145 : data_rom <= {16'd30098, 16'd12953};
                15'd12146 : data_rom <= {16'd30100, 16'd12950};
                15'd12147 : data_rom <= {16'd30101, 16'd12947};
                15'd12148 : data_rom <= {16'd30102, 16'd12945};
                15'd12149 : data_rom <= {16'd30103, 16'd12942};
                15'd12150 : data_rom <= {16'd30105, 16'd12939};
                15'd12151 : data_rom <= {16'd30106, 16'd12936};
                15'd12152 : data_rom <= {16'd30107, 16'd12933};
                15'd12153 : data_rom <= {16'd30108, 16'd12930};
                15'd12154 : data_rom <= {16'd30110, 16'd12927};
                15'd12155 : data_rom <= {16'd30111, 16'd12924};
                15'd12156 : data_rom <= {16'd30112, 16'd12921};
                15'd12157 : data_rom <= {16'd30113, 16'd12919};
                15'd12158 : data_rom <= {16'd30115, 16'd12916};
                15'd12159 : data_rom <= {16'd30116, 16'd12913};
                15'd12160 : data_rom <= {16'd30117, 16'd12910};
                15'd12161 : data_rom <= {16'd30118, 16'd12907};
                15'd12162 : data_rom <= {16'd30119, 16'd12904};
                15'd12163 : data_rom <= {16'd30121, 16'd12901};
                15'd12164 : data_rom <= {16'd30122, 16'd12898};
                15'd12165 : data_rom <= {16'd30123, 16'd12895};
                15'd12166 : data_rom <= {16'd30124, 16'd12893};
                15'd12167 : data_rom <= {16'd30126, 16'd12890};
                15'd12168 : data_rom <= {16'd30127, 16'd12887};
                15'd12169 : data_rom <= {16'd30128, 16'd12884};
                15'd12170 : data_rom <= {16'd30129, 16'd12881};
                15'd12171 : data_rom <= {16'd30131, 16'd12878};
                15'd12172 : data_rom <= {16'd30132, 16'd12875};
                15'd12173 : data_rom <= {16'd30133, 16'd12872};
                15'd12174 : data_rom <= {16'd30134, 16'd12869};
                15'd12175 : data_rom <= {16'd30136, 16'd12867};
                15'd12176 : data_rom <= {16'd30137, 16'd12864};
                15'd12177 : data_rom <= {16'd30138, 16'd12861};
                15'd12178 : data_rom <= {16'd30139, 16'd12858};
                15'd12179 : data_rom <= {16'd30140, 16'd12855};
                15'd12180 : data_rom <= {16'd30142, 16'd12852};
                15'd12181 : data_rom <= {16'd30143, 16'd12849};
                15'd12182 : data_rom <= {16'd30144, 16'd12846};
                15'd12183 : data_rom <= {16'd30145, 16'd12843};
                15'd12184 : data_rom <= {16'd30147, 16'd12841};
                15'd12185 : data_rom <= {16'd30148, 16'd12838};
                15'd12186 : data_rom <= {16'd30149, 16'd12835};
                15'd12187 : data_rom <= {16'd30150, 16'd12832};
                15'd12188 : data_rom <= {16'd30152, 16'd12829};
                15'd12189 : data_rom <= {16'd30153, 16'd12826};
                15'd12190 : data_rom <= {16'd30154, 16'd12823};
                15'd12191 : data_rom <= {16'd30155, 16'd12820};
                15'd12192 : data_rom <= {16'd30156, 16'd12817};
                15'd12193 : data_rom <= {16'd30158, 16'd12815};
                15'd12194 : data_rom <= {16'd30159, 16'd12812};
                15'd12195 : data_rom <= {16'd30160, 16'd12809};
                15'd12196 : data_rom <= {16'd30161, 16'd12806};
                15'd12197 : data_rom <= {16'd30163, 16'd12803};
                15'd12198 : data_rom <= {16'd30164, 16'd12800};
                15'd12199 : data_rom <= {16'd30165, 16'd12797};
                15'd12200 : data_rom <= {16'd30166, 16'd12794};
                15'd12201 : data_rom <= {16'd30168, 16'd12791};
                15'd12202 : data_rom <= {16'd30169, 16'd12788};
                15'd12203 : data_rom <= {16'd30170, 16'd12786};
                15'd12204 : data_rom <= {16'd30171, 16'd12783};
                15'd12205 : data_rom <= {16'd30172, 16'd12780};
                15'd12206 : data_rom <= {16'd30174, 16'd12777};
                15'd12207 : data_rom <= {16'd30175, 16'd12774};
                15'd12208 : data_rom <= {16'd30176, 16'd12771};
                15'd12209 : data_rom <= {16'd30177, 16'd12768};
                15'd12210 : data_rom <= {16'd30179, 16'd12765};
                15'd12211 : data_rom <= {16'd30180, 16'd12762};
                15'd12212 : data_rom <= {16'd30181, 16'd12760};
                15'd12213 : data_rom <= {16'd30182, 16'd12757};
                15'd12214 : data_rom <= {16'd30183, 16'd12754};
                15'd12215 : data_rom <= {16'd30185, 16'd12751};
                15'd12216 : data_rom <= {16'd30186, 16'd12748};
                15'd12217 : data_rom <= {16'd30187, 16'd12745};
                15'd12218 : data_rom <= {16'd30188, 16'd12742};
                15'd12219 : data_rom <= {16'd30190, 16'd12739};
                15'd12220 : data_rom <= {16'd30191, 16'd12736};
                15'd12221 : data_rom <= {16'd30192, 16'd12734};
                15'd12222 : data_rom <= {16'd30193, 16'd12731};
                15'd12223 : data_rom <= {16'd30194, 16'd12728};
                15'd12224 : data_rom <= {16'd30196, 16'd12725};
                15'd12225 : data_rom <= {16'd30197, 16'd12722};
                15'd12226 : data_rom <= {16'd30198, 16'd12719};
                15'd12227 : data_rom <= {16'd30199, 16'd12716};
                15'd12228 : data_rom <= {16'd30201, 16'd12713};
                15'd12229 : data_rom <= {16'd30202, 16'd12710};
                15'd12230 : data_rom <= {16'd30203, 16'd12707};
                15'd12231 : data_rom <= {16'd30204, 16'd12705};
                15'd12232 : data_rom <= {16'd30205, 16'd12702};
                15'd12233 : data_rom <= {16'd30207, 16'd12699};
                15'd12234 : data_rom <= {16'd30208, 16'd12696};
                15'd12235 : data_rom <= {16'd30209, 16'd12693};
                15'd12236 : data_rom <= {16'd30210, 16'd12690};
                15'd12237 : data_rom <= {16'd30211, 16'd12687};
                15'd12238 : data_rom <= {16'd30213, 16'd12684};
                15'd12239 : data_rom <= {16'd30214, 16'd12681};
                15'd12240 : data_rom <= {16'd30215, 16'd12678};
                15'd12241 : data_rom <= {16'd30216, 16'd12676};
                15'd12242 : data_rom <= {16'd30218, 16'd12673};
                15'd12243 : data_rom <= {16'd30219, 16'd12670};
                15'd12244 : data_rom <= {16'd30220, 16'd12667};
                15'd12245 : data_rom <= {16'd30221, 16'd12664};
                15'd12246 : data_rom <= {16'd30222, 16'd12661};
                15'd12247 : data_rom <= {16'd30224, 16'd12658};
                15'd12248 : data_rom <= {16'd30225, 16'd12655};
                15'd12249 : data_rom <= {16'd30226, 16'd12652};
                15'd12250 : data_rom <= {16'd30227, 16'd12650};
                15'd12251 : data_rom <= {16'd30228, 16'd12647};
                15'd12252 : data_rom <= {16'd30230, 16'd12644};
                15'd12253 : data_rom <= {16'd30231, 16'd12641};
                15'd12254 : data_rom <= {16'd30232, 16'd12638};
                15'd12255 : data_rom <= {16'd30233, 16'd12635};
                15'd12256 : data_rom <= {16'd30235, 16'd12632};
                15'd12257 : data_rom <= {16'd30236, 16'd12629};
                15'd12258 : data_rom <= {16'd30237, 16'd12626};
                15'd12259 : data_rom <= {16'd30238, 16'd12623};
                15'd12260 : data_rom <= {16'd30239, 16'd12621};
                15'd12261 : data_rom <= {16'd30241, 16'd12618};
                15'd12262 : data_rom <= {16'd30242, 16'd12615};
                15'd12263 : data_rom <= {16'd30243, 16'd12612};
                15'd12264 : data_rom <= {16'd30244, 16'd12609};
                15'd12265 : data_rom <= {16'd30245, 16'd12606};
                15'd12266 : data_rom <= {16'd30247, 16'd12603};
                15'd12267 : data_rom <= {16'd30248, 16'd12600};
                15'd12268 : data_rom <= {16'd30249, 16'd12597};
                15'd12269 : data_rom <= {16'd30250, 16'd12594};
                15'd12270 : data_rom <= {16'd30251, 16'd12592};
                15'd12271 : data_rom <= {16'd30253, 16'd12589};
                15'd12272 : data_rom <= {16'd30254, 16'd12586};
                15'd12273 : data_rom <= {16'd30255, 16'd12583};
                15'd12274 : data_rom <= {16'd30256, 16'd12580};
                15'd12275 : data_rom <= {16'd30258, 16'd12577};
                15'd12276 : data_rom <= {16'd30259, 16'd12574};
                15'd12277 : data_rom <= {16'd30260, 16'd12571};
                15'd12278 : data_rom <= {16'd30261, 16'd12568};
                15'd12279 : data_rom <= {16'd30262, 16'd12565};
                15'd12280 : data_rom <= {16'd30264, 16'd12563};
                15'd12281 : data_rom <= {16'd30265, 16'd12560};
                15'd12282 : data_rom <= {16'd30266, 16'd12557};
                15'd12283 : data_rom <= {16'd30267, 16'd12554};
                15'd12284 : data_rom <= {16'd30268, 16'd12551};
                15'd12285 : data_rom <= {16'd30270, 16'd12548};
                15'd12286 : data_rom <= {16'd30271, 16'd12545};
                15'd12287 : data_rom <= {16'd30272, 16'd12542};
                15'd12288 : data_rom <= {16'd30273, 16'd12539};
                15'd12289 : data_rom <= {16'd30274, 16'd12536};
                15'd12290 : data_rom <= {16'd30276, 16'd12533};
                15'd12291 : data_rom <= {16'd30277, 16'd12531};
                15'd12292 : data_rom <= {16'd30278, 16'd12528};
                15'd12293 : data_rom <= {16'd30279, 16'd12525};
                15'd12294 : data_rom <= {16'd30280, 16'd12522};
                15'd12295 : data_rom <= {16'd30282, 16'd12519};
                15'd12296 : data_rom <= {16'd30283, 16'd12516};
                15'd12297 : data_rom <= {16'd30284, 16'd12513};
                15'd12298 : data_rom <= {16'd30285, 16'd12510};
                15'd12299 : data_rom <= {16'd30286, 16'd12507};
                15'd12300 : data_rom <= {16'd30288, 16'd12504};
                15'd12301 : data_rom <= {16'd30289, 16'd12502};
                15'd12302 : data_rom <= {16'd30290, 16'd12499};
                15'd12303 : data_rom <= {16'd30291, 16'd12496};
                15'd12304 : data_rom <= {16'd30292, 16'd12493};
                15'd12305 : data_rom <= {16'd30294, 16'd12490};
                15'd12306 : data_rom <= {16'd30295, 16'd12487};
                15'd12307 : data_rom <= {16'd30296, 16'd12484};
                15'd12308 : data_rom <= {16'd30297, 16'd12481};
                15'd12309 : data_rom <= {16'd30298, 16'd12478};
                15'd12310 : data_rom <= {16'd30300, 16'd12475};
                15'd12311 : data_rom <= {16'd30301, 16'd12473};
                15'd12312 : data_rom <= {16'd30302, 16'd12470};
                15'd12313 : data_rom <= {16'd30303, 16'd12467};
                15'd12314 : data_rom <= {16'd30304, 16'd12464};
                15'd12315 : data_rom <= {16'd30306, 16'd12461};
                15'd12316 : data_rom <= {16'd30307, 16'd12458};
                15'd12317 : data_rom <= {16'd30308, 16'd12455};
                15'd12318 : data_rom <= {16'd30309, 16'd12452};
                15'd12319 : data_rom <= {16'd30310, 16'd12449};
                15'd12320 : data_rom <= {16'd30311, 16'd12446};
                15'd12321 : data_rom <= {16'd30313, 16'd12443};
                15'd12322 : data_rom <= {16'd30314, 16'd12441};
                15'd12323 : data_rom <= {16'd30315, 16'd12438};
                15'd12324 : data_rom <= {16'd30316, 16'd12435};
                15'd12325 : data_rom <= {16'd30317, 16'd12432};
                15'd12326 : data_rom <= {16'd30319, 16'd12429};
                15'd12327 : data_rom <= {16'd30320, 16'd12426};
                15'd12328 : data_rom <= {16'd30321, 16'd12423};
                15'd12329 : data_rom <= {16'd30322, 16'd12420};
                15'd12330 : data_rom <= {16'd30323, 16'd12417};
                15'd12331 : data_rom <= {16'd30325, 16'd12414};
                15'd12332 : data_rom <= {16'd30326, 16'd12411};
                15'd12333 : data_rom <= {16'd30327, 16'd12409};
                15'd12334 : data_rom <= {16'd30328, 16'd12406};
                15'd12335 : data_rom <= {16'd30329, 16'd12403};
                15'd12336 : data_rom <= {16'd30331, 16'd12400};
                15'd12337 : data_rom <= {16'd30332, 16'd12397};
                15'd12338 : data_rom <= {16'd30333, 16'd12394};
                15'd12339 : data_rom <= {16'd30334, 16'd12391};
                15'd12340 : data_rom <= {16'd30335, 16'd12388};
                15'd12341 : data_rom <= {16'd30336, 16'd12385};
                15'd12342 : data_rom <= {16'd30338, 16'd12382};
                15'd12343 : data_rom <= {16'd30339, 16'd12379};
                15'd12344 : data_rom <= {16'd30340, 16'd12377};
                15'd12345 : data_rom <= {16'd30341, 16'd12374};
                15'd12346 : data_rom <= {16'd30342, 16'd12371};
                15'd12347 : data_rom <= {16'd30344, 16'd12368};
                15'd12348 : data_rom <= {16'd30345, 16'd12365};
                15'd12349 : data_rom <= {16'd30346, 16'd12362};
                15'd12350 : data_rom <= {16'd30347, 16'd12359};
                15'd12351 : data_rom <= {16'd30348, 16'd12356};
                15'd12352 : data_rom <= {16'd30350, 16'd12353};
                15'd12353 : data_rom <= {16'd30351, 16'd12350};
                15'd12354 : data_rom <= {16'd30352, 16'd12347};
                15'd12355 : data_rom <= {16'd30353, 16'd12345};
                15'd12356 : data_rom <= {16'd30354, 16'd12342};
                15'd12357 : data_rom <= {16'd30355, 16'd12339};
                15'd12358 : data_rom <= {16'd30357, 16'd12336};
                15'd12359 : data_rom <= {16'd30358, 16'd12333};
                15'd12360 : data_rom <= {16'd30359, 16'd12330};
                15'd12361 : data_rom <= {16'd30360, 16'd12327};
                15'd12362 : data_rom <= {16'd30361, 16'd12324};
                15'd12363 : data_rom <= {16'd30363, 16'd12321};
                15'd12364 : data_rom <= {16'd30364, 16'd12318};
                15'd12365 : data_rom <= {16'd30365, 16'd12315};
                15'd12366 : data_rom <= {16'd30366, 16'd12313};
                15'd12367 : data_rom <= {16'd30367, 16'd12310};
                15'd12368 : data_rom <= {16'd30368, 16'd12307};
                15'd12369 : data_rom <= {16'd30370, 16'd12304};
                15'd12370 : data_rom <= {16'd30371, 16'd12301};
                15'd12371 : data_rom <= {16'd30372, 16'd12298};
                15'd12372 : data_rom <= {16'd30373, 16'd12295};
                15'd12373 : data_rom <= {16'd30374, 16'd12292};
                15'd12374 : data_rom <= {16'd30376, 16'd12289};
                15'd12375 : data_rom <= {16'd30377, 16'd12286};
                15'd12376 : data_rom <= {16'd30378, 16'd12283};
                15'd12377 : data_rom <= {16'd30379, 16'd12281};
                15'd12378 : data_rom <= {16'd30380, 16'd12278};
                15'd12379 : data_rom <= {16'd30381, 16'd12275};
                15'd12380 : data_rom <= {16'd30383, 16'd12272};
                15'd12381 : data_rom <= {16'd30384, 16'd12269};
                15'd12382 : data_rom <= {16'd30385, 16'd12266};
                15'd12383 : data_rom <= {16'd30386, 16'd12263};
                15'd12384 : data_rom <= {16'd30387, 16'd12260};
                15'd12385 : data_rom <= {16'd30388, 16'd12257};
                15'd12386 : data_rom <= {16'd30390, 16'd12254};
                15'd12387 : data_rom <= {16'd30391, 16'd12251};
                15'd12388 : data_rom <= {16'd30392, 16'd12248};
                15'd12389 : data_rom <= {16'd30393, 16'd12246};
                15'd12390 : data_rom <= {16'd30394, 16'd12243};
                15'd12391 : data_rom <= {16'd30396, 16'd12240};
                15'd12392 : data_rom <= {16'd30397, 16'd12237};
                15'd12393 : data_rom <= {16'd30398, 16'd12234};
                15'd12394 : data_rom <= {16'd30399, 16'd12231};
                15'd12395 : data_rom <= {16'd30400, 16'd12228};
                15'd12396 : data_rom <= {16'd30401, 16'd12225};
                15'd12397 : data_rom <= {16'd30403, 16'd12222};
                15'd12398 : data_rom <= {16'd30404, 16'd12219};
                15'd12399 : data_rom <= {16'd30405, 16'd12216};
                15'd12400 : data_rom <= {16'd30406, 16'd12214};
                15'd12401 : data_rom <= {16'd30407, 16'd12211};
                15'd12402 : data_rom <= {16'd30408, 16'd12208};
                15'd12403 : data_rom <= {16'd30410, 16'd12205};
                15'd12404 : data_rom <= {16'd30411, 16'd12202};
                15'd12405 : data_rom <= {16'd30412, 16'd12199};
                15'd12406 : data_rom <= {16'd30413, 16'd12196};
                15'd12407 : data_rom <= {16'd30414, 16'd12193};
                15'd12408 : data_rom <= {16'd30415, 16'd12190};
                15'd12409 : data_rom <= {16'd30417, 16'd12187};
                15'd12410 : data_rom <= {16'd30418, 16'd12184};
                15'd12411 : data_rom <= {16'd30419, 16'd12181};
                15'd12412 : data_rom <= {16'd30420, 16'd12179};
                15'd12413 : data_rom <= {16'd30421, 16'd12176};
                15'd12414 : data_rom <= {16'd30422, 16'd12173};
                15'd12415 : data_rom <= {16'd30424, 16'd12170};
                15'd12416 : data_rom <= {16'd30425, 16'd12167};
                15'd12417 : data_rom <= {16'd30426, 16'd12164};
                15'd12418 : data_rom <= {16'd30427, 16'd12161};
                15'd12419 : data_rom <= {16'd30428, 16'd12158};
                15'd12420 : data_rom <= {16'd30429, 16'd12155};
                15'd12421 : data_rom <= {16'd30431, 16'd12152};
                15'd12422 : data_rom <= {16'd30432, 16'd12149};
                15'd12423 : data_rom <= {16'd30433, 16'd12146};
                15'd12424 : data_rom <= {16'd30434, 16'd12144};
                15'd12425 : data_rom <= {16'd30435, 16'd12141};
                15'd12426 : data_rom <= {16'd30436, 16'd12138};
                15'd12427 : data_rom <= {16'd30438, 16'd12135};
                15'd12428 : data_rom <= {16'd30439, 16'd12132};
                15'd12429 : data_rom <= {16'd30440, 16'd12129};
                15'd12430 : data_rom <= {16'd30441, 16'd12126};
                15'd12431 : data_rom <= {16'd30442, 16'd12123};
                15'd12432 : data_rom <= {16'd30443, 16'd12120};
                15'd12433 : data_rom <= {16'd30445, 16'd12117};
                15'd12434 : data_rom <= {16'd30446, 16'd12114};
                15'd12435 : data_rom <= {16'd30447, 16'd12111};
                15'd12436 : data_rom <= {16'd30448, 16'd12108};
                15'd12437 : data_rom <= {16'd30449, 16'd12106};
                15'd12438 : data_rom <= {16'd30450, 16'd12103};
                15'd12439 : data_rom <= {16'd30452, 16'd12100};
                15'd12440 : data_rom <= {16'd30453, 16'd12097};
                15'd12441 : data_rom <= {16'd30454, 16'd12094};
                15'd12442 : data_rom <= {16'd30455, 16'd12091};
                15'd12443 : data_rom <= {16'd30456, 16'd12088};
                15'd12444 : data_rom <= {16'd30457, 16'd12085};
                15'd12445 : data_rom <= {16'd30458, 16'd12082};
                15'd12446 : data_rom <= {16'd30460, 16'd12079};
                15'd12447 : data_rom <= {16'd30461, 16'd12076};
                15'd12448 : data_rom <= {16'd30462, 16'd12073};
                15'd12449 : data_rom <= {16'd30463, 16'd12071};
                15'd12450 : data_rom <= {16'd30464, 16'd12068};
                15'd12451 : data_rom <= {16'd30465, 16'd12065};
                15'd12452 : data_rom <= {16'd30467, 16'd12062};
                15'd12453 : data_rom <= {16'd30468, 16'd12059};
                15'd12454 : data_rom <= {16'd30469, 16'd12056};
                15'd12455 : data_rom <= {16'd30470, 16'd12053};
                15'd12456 : data_rom <= {16'd30471, 16'd12050};
                15'd12457 : data_rom <= {16'd30472, 16'd12047};
                15'd12458 : data_rom <= {16'd30474, 16'd12044};
                15'd12459 : data_rom <= {16'd30475, 16'd12041};
                15'd12460 : data_rom <= {16'd30476, 16'd12038};
                15'd12461 : data_rom <= {16'd30477, 16'd12035};
                15'd12462 : data_rom <= {16'd30478, 16'd12033};
                15'd12463 : data_rom <= {16'd30479, 16'd12030};
                15'd12464 : data_rom <= {16'd30480, 16'd12027};
                15'd12465 : data_rom <= {16'd30482, 16'd12024};
                15'd12466 : data_rom <= {16'd30483, 16'd12021};
                15'd12467 : data_rom <= {16'd30484, 16'd12018};
                15'd12468 : data_rom <= {16'd30485, 16'd12015};
                15'd12469 : data_rom <= {16'd30486, 16'd12012};
                15'd12470 : data_rom <= {16'd30487, 16'd12009};
                15'd12471 : data_rom <= {16'd30489, 16'd12006};
                15'd12472 : data_rom <= {16'd30490, 16'd12003};
                15'd12473 : data_rom <= {16'd30491, 16'd12000};
                15'd12474 : data_rom <= {16'd30492, 16'd11997};
                15'd12475 : data_rom <= {16'd30493, 16'd11995};
                15'd12476 : data_rom <= {16'd30494, 16'd11992};
                15'd12477 : data_rom <= {16'd30495, 16'd11989};
                15'd12478 : data_rom <= {16'd30497, 16'd11986};
                15'd12479 : data_rom <= {16'd30498, 16'd11983};
                15'd12480 : data_rom <= {16'd30499, 16'd11980};
                15'd12481 : data_rom <= {16'd30500, 16'd11977};
                15'd12482 : data_rom <= {16'd30501, 16'd11974};
                15'd12483 : data_rom <= {16'd30502, 16'd11971};
                15'd12484 : data_rom <= {16'd30503, 16'd11968};
                15'd12485 : data_rom <= {16'd30505, 16'd11965};
                15'd12486 : data_rom <= {16'd30506, 16'd11962};
                15'd12487 : data_rom <= {16'd30507, 16'd11959};
                15'd12488 : data_rom <= {16'd30508, 16'd11957};
                15'd12489 : data_rom <= {16'd30509, 16'd11954};
                15'd12490 : data_rom <= {16'd30510, 16'd11951};
                15'd12491 : data_rom <= {16'd30511, 16'd11948};
                15'd12492 : data_rom <= {16'd30513, 16'd11945};
                15'd12493 : data_rom <= {16'd30514, 16'd11942};
                15'd12494 : data_rom <= {16'd30515, 16'd11939};
                15'd12495 : data_rom <= {16'd30516, 16'd11936};
                15'd12496 : data_rom <= {16'd30517, 16'd11933};
                15'd12497 : data_rom <= {16'd30518, 16'd11930};
                15'd12498 : data_rom <= {16'd30519, 16'd11927};
                15'd12499 : data_rom <= {16'd30521, 16'd11924};
                15'd12500 : data_rom <= {16'd30522, 16'd11921};
                15'd12501 : data_rom <= {16'd30523, 16'd11919};
                15'd12502 : data_rom <= {16'd30524, 16'd11916};
                15'd12503 : data_rom <= {16'd30525, 16'd11913};
                15'd12504 : data_rom <= {16'd30526, 16'd11910};
                15'd12505 : data_rom <= {16'd30527, 16'd11907};
                15'd12506 : data_rom <= {16'd30529, 16'd11904};
                15'd12507 : data_rom <= {16'd30530, 16'd11901};
                15'd12508 : data_rom <= {16'd30531, 16'd11898};
                15'd12509 : data_rom <= {16'd30532, 16'd11895};
                15'd12510 : data_rom <= {16'd30533, 16'd11892};
                15'd12511 : data_rom <= {16'd30534, 16'd11889};
                15'd12512 : data_rom <= {16'd30535, 16'd11886};
                15'd12513 : data_rom <= {16'd30537, 16'd11883};
                15'd12514 : data_rom <= {16'd30538, 16'd11880};
                15'd12515 : data_rom <= {16'd30539, 16'd11878};
                15'd12516 : data_rom <= {16'd30540, 16'd11875};
                15'd12517 : data_rom <= {16'd30541, 16'd11872};
                15'd12518 : data_rom <= {16'd30542, 16'd11869};
                15'd12519 : data_rom <= {16'd30543, 16'd11866};
                15'd12520 : data_rom <= {16'd30545, 16'd11863};
                15'd12521 : data_rom <= {16'd30546, 16'd11860};
                15'd12522 : data_rom <= {16'd30547, 16'd11857};
                15'd12523 : data_rom <= {16'd30548, 16'd11854};
                15'd12524 : data_rom <= {16'd30549, 16'd11851};
                15'd12525 : data_rom <= {16'd30550, 16'd11848};
                15'd12526 : data_rom <= {16'd30551, 16'd11845};
                15'd12527 : data_rom <= {16'd30553, 16'd11842};
                15'd12528 : data_rom <= {16'd30554, 16'd11839};
                15'd12529 : data_rom <= {16'd30555, 16'd11837};
                15'd12530 : data_rom <= {16'd30556, 16'd11834};
                15'd12531 : data_rom <= {16'd30557, 16'd11831};
                15'd12532 : data_rom <= {16'd30558, 16'd11828};
                15'd12533 : data_rom <= {16'd30559, 16'd11825};
                15'd12534 : data_rom <= {16'd30560, 16'd11822};
                15'd12535 : data_rom <= {16'd30562, 16'd11819};
                15'd12536 : data_rom <= {16'd30563, 16'd11816};
                15'd12537 : data_rom <= {16'd30564, 16'd11813};
                15'd12538 : data_rom <= {16'd30565, 16'd11810};
                15'd12539 : data_rom <= {16'd30566, 16'd11807};
                15'd12540 : data_rom <= {16'd30567, 16'd11804};
                15'd12541 : data_rom <= {16'd30568, 16'd11801};
                15'd12542 : data_rom <= {16'd30570, 16'd11798};
                15'd12543 : data_rom <= {16'd30571, 16'd11796};
                15'd12544 : data_rom <= {16'd30572, 16'd11793};
                15'd12545 : data_rom <= {16'd30573, 16'd11790};
                15'd12546 : data_rom <= {16'd30574, 16'd11787};
                15'd12547 : data_rom <= {16'd30575, 16'd11784};
                15'd12548 : data_rom <= {16'd30576, 16'd11781};
                15'd12549 : data_rom <= {16'd30577, 16'd11778};
                15'd12550 : data_rom <= {16'd30579, 16'd11775};
                15'd12551 : data_rom <= {16'd30580, 16'd11772};
                15'd12552 : data_rom <= {16'd30581, 16'd11769};
                15'd12553 : data_rom <= {16'd30582, 16'd11766};
                15'd12554 : data_rom <= {16'd30583, 16'd11763};
                15'd12555 : data_rom <= {16'd30584, 16'd11760};
                15'd12556 : data_rom <= {16'd30585, 16'd11757};
                15'd12557 : data_rom <= {16'd30586, 16'd11754};
                15'd12558 : data_rom <= {16'd30588, 16'd11752};
                15'd12559 : data_rom <= {16'd30589, 16'd11749};
                15'd12560 : data_rom <= {16'd30590, 16'd11746};
                15'd12561 : data_rom <= {16'd30591, 16'd11743};
                15'd12562 : data_rom <= {16'd30592, 16'd11740};
                15'd12563 : data_rom <= {16'd30593, 16'd11737};
                15'd12564 : data_rom <= {16'd30594, 16'd11734};
                15'd12565 : data_rom <= {16'd30595, 16'd11731};
                15'd12566 : data_rom <= {16'd30597, 16'd11728};
                15'd12567 : data_rom <= {16'd30598, 16'd11725};
                15'd12568 : data_rom <= {16'd30599, 16'd11722};
                15'd12569 : data_rom <= {16'd30600, 16'd11719};
                15'd12570 : data_rom <= {16'd30601, 16'd11716};
                15'd12571 : data_rom <= {16'd30602, 16'd11713};
                15'd12572 : data_rom <= {16'd30603, 16'd11710};
                15'd12573 : data_rom <= {16'd30604, 16'd11708};
                15'd12574 : data_rom <= {16'd30606, 16'd11705};
                15'd12575 : data_rom <= {16'd30607, 16'd11702};
                15'd12576 : data_rom <= {16'd30608, 16'd11699};
                15'd12577 : data_rom <= {16'd30609, 16'd11696};
                15'd12578 : data_rom <= {16'd30610, 16'd11693};
                15'd12579 : data_rom <= {16'd30611, 16'd11690};
                15'd12580 : data_rom <= {16'd30612, 16'd11687};
                15'd12581 : data_rom <= {16'd30613, 16'd11684};
                15'd12582 : data_rom <= {16'd30615, 16'd11681};
                15'd12583 : data_rom <= {16'd30616, 16'd11678};
                15'd12584 : data_rom <= {16'd30617, 16'd11675};
                15'd12585 : data_rom <= {16'd30618, 16'd11672};
                15'd12586 : data_rom <= {16'd30619, 16'd11669};
                15'd12587 : data_rom <= {16'd30620, 16'd11666};
                15'd12588 : data_rom <= {16'd30621, 16'd11664};
                15'd12589 : data_rom <= {16'd30622, 16'd11661};
                15'd12590 : data_rom <= {16'd30624, 16'd11658};
                15'd12591 : data_rom <= {16'd30625, 16'd11655};
                15'd12592 : data_rom <= {16'd30626, 16'd11652};
                15'd12593 : data_rom <= {16'd30627, 16'd11649};
                15'd12594 : data_rom <= {16'd30628, 16'd11646};
                15'd12595 : data_rom <= {16'd30629, 16'd11643};
                15'd12596 : data_rom <= {16'd30630, 16'd11640};
                15'd12597 : data_rom <= {16'd30631, 16'd11637};
                15'd12598 : data_rom <= {16'd30632, 16'd11634};
                15'd12599 : data_rom <= {16'd30634, 16'd11631};
                15'd12600 : data_rom <= {16'd30635, 16'd11628};
                15'd12601 : data_rom <= {16'd30636, 16'd11625};
                15'd12602 : data_rom <= {16'd30637, 16'd11622};
                15'd12603 : data_rom <= {16'd30638, 16'd11619};
                15'd12604 : data_rom <= {16'd30639, 16'd11617};
                15'd12605 : data_rom <= {16'd30640, 16'd11614};
                15'd12606 : data_rom <= {16'd30641, 16'd11611};
                15'd12607 : data_rom <= {16'd30642, 16'd11608};
                15'd12608 : data_rom <= {16'd30644, 16'd11605};
                15'd12609 : data_rom <= {16'd30645, 16'd11602};
                15'd12610 : data_rom <= {16'd30646, 16'd11599};
                15'd12611 : data_rom <= {16'd30647, 16'd11596};
                15'd12612 : data_rom <= {16'd30648, 16'd11593};
                15'd12613 : data_rom <= {16'd30649, 16'd11590};
                15'd12614 : data_rom <= {16'd30650, 16'd11587};
                15'd12615 : data_rom <= {16'd30651, 16'd11584};
                15'd12616 : data_rom <= {16'd30652, 16'd11581};
                15'd12617 : data_rom <= {16'd30654, 16'd11578};
                15'd12618 : data_rom <= {16'd30655, 16'd11575};
                15'd12619 : data_rom <= {16'd30656, 16'd11572};
                15'd12620 : data_rom <= {16'd30657, 16'd11570};
                15'd12621 : data_rom <= {16'd30658, 16'd11567};
                15'd12622 : data_rom <= {16'd30659, 16'd11564};
                15'd12623 : data_rom <= {16'd30660, 16'd11561};
                15'd12624 : data_rom <= {16'd30661, 16'd11558};
                15'd12625 : data_rom <= {16'd30662, 16'd11555};
                15'd12626 : data_rom <= {16'd30664, 16'd11552};
                15'd12627 : data_rom <= {16'd30665, 16'd11549};
                15'd12628 : data_rom <= {16'd30666, 16'd11546};
                15'd12629 : data_rom <= {16'd30667, 16'd11543};
                15'd12630 : data_rom <= {16'd30668, 16'd11540};
                15'd12631 : data_rom <= {16'd30669, 16'd11537};
                15'd12632 : data_rom <= {16'd30670, 16'd11534};
                15'd12633 : data_rom <= {16'd30671, 16'd11531};
                15'd12634 : data_rom <= {16'd30672, 16'd11528};
                15'd12635 : data_rom <= {16'd30674, 16'd11525};
                15'd12636 : data_rom <= {16'd30675, 16'd11522};
                15'd12637 : data_rom <= {16'd30676, 16'd11520};
                15'd12638 : data_rom <= {16'd30677, 16'd11517};
                15'd12639 : data_rom <= {16'd30678, 16'd11514};
                15'd12640 : data_rom <= {16'd30679, 16'd11511};
                15'd12641 : data_rom <= {16'd30680, 16'd11508};
                15'd12642 : data_rom <= {16'd30681, 16'd11505};
                15'd12643 : data_rom <= {16'd30682, 16'd11502};
                15'd12644 : data_rom <= {16'd30683, 16'd11499};
                15'd12645 : data_rom <= {16'd30685, 16'd11496};
                15'd12646 : data_rom <= {16'd30686, 16'd11493};
                15'd12647 : data_rom <= {16'd30687, 16'd11490};
                15'd12648 : data_rom <= {16'd30688, 16'd11487};
                15'd12649 : data_rom <= {16'd30689, 16'd11484};
                15'd12650 : data_rom <= {16'd30690, 16'd11481};
                15'd12651 : data_rom <= {16'd30691, 16'd11478};
                15'd12652 : data_rom <= {16'd30692, 16'd11475};
                15'd12653 : data_rom <= {16'd30693, 16'd11472};
                15'd12654 : data_rom <= {16'd30694, 16'd11470};
                15'd12655 : data_rom <= {16'd30696, 16'd11467};
                15'd12656 : data_rom <= {16'd30697, 16'd11464};
                15'd12657 : data_rom <= {16'd30698, 16'd11461};
                15'd12658 : data_rom <= {16'd30699, 16'd11458};
                15'd12659 : data_rom <= {16'd30700, 16'd11455};
                15'd12660 : data_rom <= {16'd30701, 16'd11452};
                15'd12661 : data_rom <= {16'd30702, 16'd11449};
                15'd12662 : data_rom <= {16'd30703, 16'd11446};
                15'd12663 : data_rom <= {16'd30704, 16'd11443};
                15'd12664 : data_rom <= {16'd30705, 16'd11440};
                15'd12665 : data_rom <= {16'd30707, 16'd11437};
                15'd12666 : data_rom <= {16'd30708, 16'd11434};
                15'd12667 : data_rom <= {16'd30709, 16'd11431};
                15'd12668 : data_rom <= {16'd30710, 16'd11428};
                15'd12669 : data_rom <= {16'd30711, 16'd11425};
                15'd12670 : data_rom <= {16'd30712, 16'd11422};
                15'd12671 : data_rom <= {16'd30713, 16'd11419};
                15'd12672 : data_rom <= {16'd30714, 16'd11417};
                15'd12673 : data_rom <= {16'd30715, 16'd11414};
                15'd12674 : data_rom <= {16'd30716, 16'd11411};
                15'd12675 : data_rom <= {16'd30717, 16'd11408};
                15'd12676 : data_rom <= {16'd30719, 16'd11405};
                15'd12677 : data_rom <= {16'd30720, 16'd11402};
                15'd12678 : data_rom <= {16'd30721, 16'd11399};
                15'd12679 : data_rom <= {16'd30722, 16'd11396};
                15'd12680 : data_rom <= {16'd30723, 16'd11393};
                15'd12681 : data_rom <= {16'd30724, 16'd11390};
                15'd12682 : data_rom <= {16'd30725, 16'd11387};
                15'd12683 : data_rom <= {16'd30726, 16'd11384};
                15'd12684 : data_rom <= {16'd30727, 16'd11381};
                15'd12685 : data_rom <= {16'd30728, 16'd11378};
                15'd12686 : data_rom <= {16'd30730, 16'd11375};
                15'd12687 : data_rom <= {16'd30731, 16'd11372};
                15'd12688 : data_rom <= {16'd30732, 16'd11369};
                15'd12689 : data_rom <= {16'd30733, 16'd11366};
                15'd12690 : data_rom <= {16'd30734, 16'd11363};
                15'd12691 : data_rom <= {16'd30735, 16'd11361};
                15'd12692 : data_rom <= {16'd30736, 16'd11358};
                15'd12693 : data_rom <= {16'd30737, 16'd11355};
                15'd12694 : data_rom <= {16'd30738, 16'd11352};
                15'd12695 : data_rom <= {16'd30739, 16'd11349};
                15'd12696 : data_rom <= {16'd30740, 16'd11346};
                15'd12697 : data_rom <= {16'd30741, 16'd11343};
                15'd12698 : data_rom <= {16'd30743, 16'd11340};
                15'd12699 : data_rom <= {16'd30744, 16'd11337};
                15'd12700 : data_rom <= {16'd30745, 16'd11334};
                15'd12701 : data_rom <= {16'd30746, 16'd11331};
                15'd12702 : data_rom <= {16'd30747, 16'd11328};
                15'd12703 : data_rom <= {16'd30748, 16'd11325};
                15'd12704 : data_rom <= {16'd30749, 16'd11322};
                15'd12705 : data_rom <= {16'd30750, 16'd11319};
                15'd12706 : data_rom <= {16'd30751, 16'd11316};
                15'd12707 : data_rom <= {16'd30752, 16'd11313};
                15'd12708 : data_rom <= {16'd30753, 16'd11310};
                15'd12709 : data_rom <= {16'd30755, 16'd11307};
                15'd12710 : data_rom <= {16'd30756, 16'd11305};
                15'd12711 : data_rom <= {16'd30757, 16'd11302};
                15'd12712 : data_rom <= {16'd30758, 16'd11299};
                15'd12713 : data_rom <= {16'd30759, 16'd11296};
                15'd12714 : data_rom <= {16'd30760, 16'd11293};
                15'd12715 : data_rom <= {16'd30761, 16'd11290};
                15'd12716 : data_rom <= {16'd30762, 16'd11287};
                15'd12717 : data_rom <= {16'd30763, 16'd11284};
                15'd12718 : data_rom <= {16'd30764, 16'd11281};
                15'd12719 : data_rom <= {16'd30765, 16'd11278};
                15'd12720 : data_rom <= {16'd30766, 16'd11275};
                15'd12721 : data_rom <= {16'd30768, 16'd11272};
                15'd12722 : data_rom <= {16'd30769, 16'd11269};
                15'd12723 : data_rom <= {16'd30770, 16'd11266};
                15'd12724 : data_rom <= {16'd30771, 16'd11263};
                15'd12725 : data_rom <= {16'd30772, 16'd11260};
                15'd12726 : data_rom <= {16'd30773, 16'd11257};
                15'd12727 : data_rom <= {16'd30774, 16'd11254};
                15'd12728 : data_rom <= {16'd30775, 16'd11251};
                15'd12729 : data_rom <= {16'd30776, 16'd11248};
                15'd12730 : data_rom <= {16'd30777, 16'd11246};
                15'd12731 : data_rom <= {16'd30778, 16'd11243};
                15'd12732 : data_rom <= {16'd30779, 16'd11240};
                15'd12733 : data_rom <= {16'd30780, 16'd11237};
                15'd12734 : data_rom <= {16'd30782, 16'd11234};
                15'd12735 : data_rom <= {16'd30783, 16'd11231};
                15'd12736 : data_rom <= {16'd30784, 16'd11228};
                15'd12737 : data_rom <= {16'd30785, 16'd11225};
                15'd12738 : data_rom <= {16'd30786, 16'd11222};
                15'd12739 : data_rom <= {16'd30787, 16'd11219};
                15'd12740 : data_rom <= {16'd30788, 16'd11216};
                15'd12741 : data_rom <= {16'd30789, 16'd11213};
                15'd12742 : data_rom <= {16'd30790, 16'd11210};
                15'd12743 : data_rom <= {16'd30791, 16'd11207};
                15'd12744 : data_rom <= {16'd30792, 16'd11204};
                15'd12745 : data_rom <= {16'd30793, 16'd11201};
                15'd12746 : data_rom <= {16'd30794, 16'd11198};
                15'd12747 : data_rom <= {16'd30796, 16'd11195};
                15'd12748 : data_rom <= {16'd30797, 16'd11192};
                15'd12749 : data_rom <= {16'd30798, 16'd11189};
                15'd12750 : data_rom <= {16'd30799, 16'd11187};
                15'd12751 : data_rom <= {16'd30800, 16'd11184};
                15'd12752 : data_rom <= {16'd30801, 16'd11181};
                15'd12753 : data_rom <= {16'd30802, 16'd11178};
                15'd12754 : data_rom <= {16'd30803, 16'd11175};
                15'd12755 : data_rom <= {16'd30804, 16'd11172};
                15'd12756 : data_rom <= {16'd30805, 16'd11169};
                15'd12757 : data_rom <= {16'd30806, 16'd11166};
                15'd12758 : data_rom <= {16'd30807, 16'd11163};
                15'd12759 : data_rom <= {16'd30808, 16'd11160};
                15'd12760 : data_rom <= {16'd30809, 16'd11157};
                15'd12761 : data_rom <= {16'd30811, 16'd11154};
                15'd12762 : data_rom <= {16'd30812, 16'd11151};
                15'd12763 : data_rom <= {16'd30813, 16'd11148};
                15'd12764 : data_rom <= {16'd30814, 16'd11145};
                15'd12765 : data_rom <= {16'd30815, 16'd11142};
                15'd12766 : data_rom <= {16'd30816, 16'd11139};
                15'd12767 : data_rom <= {16'd30817, 16'd11136};
                15'd12768 : data_rom <= {16'd30818, 16'd11133};
                15'd12769 : data_rom <= {16'd30819, 16'd11130};
                15'd12770 : data_rom <= {16'd30820, 16'd11127};
                15'd12771 : data_rom <= {16'd30821, 16'd11124};
                15'd12772 : data_rom <= {16'd30822, 16'd11122};
                15'd12773 : data_rom <= {16'd30823, 16'd11119};
                15'd12774 : data_rom <= {16'd30824, 16'd11116};
                15'd12775 : data_rom <= {16'd30825, 16'd11113};
                15'd12776 : data_rom <= {16'd30827, 16'd11110};
                15'd12777 : data_rom <= {16'd30828, 16'd11107};
                15'd12778 : data_rom <= {16'd30829, 16'd11104};
                15'd12779 : data_rom <= {16'd30830, 16'd11101};
                15'd12780 : data_rom <= {16'd30831, 16'd11098};
                15'd12781 : data_rom <= {16'd30832, 16'd11095};
                15'd12782 : data_rom <= {16'd30833, 16'd11092};
                15'd12783 : data_rom <= {16'd30834, 16'd11089};
                15'd12784 : data_rom <= {16'd30835, 16'd11086};
                15'd12785 : data_rom <= {16'd30836, 16'd11083};
                15'd12786 : data_rom <= {16'd30837, 16'd11080};
                15'd12787 : data_rom <= {16'd30838, 16'd11077};
                15'd12788 : data_rom <= {16'd30839, 16'd11074};
                15'd12789 : data_rom <= {16'd30840, 16'd11071};
                15'd12790 : data_rom <= {16'd30841, 16'd11068};
                15'd12791 : data_rom <= {16'd30842, 16'd11065};
                15'd12792 : data_rom <= {16'd30844, 16'd11062};
                15'd12793 : data_rom <= {16'd30845, 16'd11059};
                15'd12794 : data_rom <= {16'd30846, 16'd11056};
                15'd12795 : data_rom <= {16'd30847, 16'd11054};
                15'd12796 : data_rom <= {16'd30848, 16'd11051};
                15'd12797 : data_rom <= {16'd30849, 16'd11048};
                15'd12798 : data_rom <= {16'd30850, 16'd11045};
                15'd12799 : data_rom <= {16'd30851, 16'd11042};
                15'd12800 : data_rom <= {16'd30852, 16'd11039};
                15'd12801 : data_rom <= {16'd30853, 16'd11036};
                15'd12802 : data_rom <= {16'd30854, 16'd11033};
                15'd12803 : data_rom <= {16'd30855, 16'd11030};
                15'd12804 : data_rom <= {16'd30856, 16'd11027};
                15'd12805 : data_rom <= {16'd30857, 16'd11024};
                15'd12806 : data_rom <= {16'd30858, 16'd11021};
                15'd12807 : data_rom <= {16'd30859, 16'd11018};
                15'd12808 : data_rom <= {16'd30860, 16'd11015};
                15'd12809 : data_rom <= {16'd30862, 16'd11012};
                15'd12810 : data_rom <= {16'd30863, 16'd11009};
                15'd12811 : data_rom <= {16'd30864, 16'd11006};
                15'd12812 : data_rom <= {16'd30865, 16'd11003};
                15'd12813 : data_rom <= {16'd30866, 16'd11000};
                15'd12814 : data_rom <= {16'd30867, 16'd10997};
                15'd12815 : data_rom <= {16'd30868, 16'd10994};
                15'd12816 : data_rom <= {16'd30869, 16'd10991};
                15'd12817 : data_rom <= {16'd30870, 16'd10988};
                15'd12818 : data_rom <= {16'd30871, 16'd10985};
                15'd12819 : data_rom <= {16'd30872, 16'd10983};
                15'd12820 : data_rom <= {16'd30873, 16'd10980};
                15'd12821 : data_rom <= {16'd30874, 16'd10977};
                15'd12822 : data_rom <= {16'd30875, 16'd10974};
                15'd12823 : data_rom <= {16'd30876, 16'd10971};
                15'd12824 : data_rom <= {16'd30877, 16'd10968};
                15'd12825 : data_rom <= {16'd30878, 16'd10965};
                15'd12826 : data_rom <= {16'd30879, 16'd10962};
                15'd12827 : data_rom <= {16'd30880, 16'd10959};
                15'd12828 : data_rom <= {16'd30882, 16'd10956};
                15'd12829 : data_rom <= {16'd30883, 16'd10953};
                15'd12830 : data_rom <= {16'd30884, 16'd10950};
                15'd12831 : data_rom <= {16'd30885, 16'd10947};
                15'd12832 : data_rom <= {16'd30886, 16'd10944};
                15'd12833 : data_rom <= {16'd30887, 16'd10941};
                15'd12834 : data_rom <= {16'd30888, 16'd10938};
                15'd12835 : data_rom <= {16'd30889, 16'd10935};
                15'd12836 : data_rom <= {16'd30890, 16'd10932};
                15'd12837 : data_rom <= {16'd30891, 16'd10929};
                15'd12838 : data_rom <= {16'd30892, 16'd10926};
                15'd12839 : data_rom <= {16'd30893, 16'd10923};
                15'd12840 : data_rom <= {16'd30894, 16'd10920};
                15'd12841 : data_rom <= {16'd30895, 16'd10917};
                15'd12842 : data_rom <= {16'd30896, 16'd10914};
                15'd12843 : data_rom <= {16'd30897, 16'd10911};
                15'd12844 : data_rom <= {16'd30898, 16'd10908};
                15'd12845 : data_rom <= {16'd30899, 16'd10906};
                15'd12846 : data_rom <= {16'd30900, 16'd10903};
                15'd12847 : data_rom <= {16'd30901, 16'd10900};
                15'd12848 : data_rom <= {16'd30902, 16'd10897};
                15'd12849 : data_rom <= {16'd30904, 16'd10894};
                15'd12850 : data_rom <= {16'd30905, 16'd10891};
                15'd12851 : data_rom <= {16'd30906, 16'd10888};
                15'd12852 : data_rom <= {16'd30907, 16'd10885};
                15'd12853 : data_rom <= {16'd30908, 16'd10882};
                15'd12854 : data_rom <= {16'd30909, 16'd10879};
                15'd12855 : data_rom <= {16'd30910, 16'd10876};
                15'd12856 : data_rom <= {16'd30911, 16'd10873};
                15'd12857 : data_rom <= {16'd30912, 16'd10870};
                15'd12858 : data_rom <= {16'd30913, 16'd10867};
                15'd12859 : data_rom <= {16'd30914, 16'd10864};
                15'd12860 : data_rom <= {16'd30915, 16'd10861};
                15'd12861 : data_rom <= {16'd30916, 16'd10858};
                15'd12862 : data_rom <= {16'd30917, 16'd10855};
                15'd12863 : data_rom <= {16'd30918, 16'd10852};
                15'd12864 : data_rom <= {16'd30919, 16'd10849};
                15'd12865 : data_rom <= {16'd30920, 16'd10846};
                15'd12866 : data_rom <= {16'd30921, 16'd10843};
                15'd12867 : data_rom <= {16'd30922, 16'd10840};
                15'd12868 : data_rom <= {16'd30923, 16'd10837};
                15'd12869 : data_rom <= {16'd30924, 16'd10834};
                15'd12870 : data_rom <= {16'd30925, 16'd10831};
                15'd12871 : data_rom <= {16'd30926, 16'd10828};
                15'd12872 : data_rom <= {16'd30927, 16'd10826};
                15'd12873 : data_rom <= {16'd30929, 16'd10823};
                15'd12874 : data_rom <= {16'd30930, 16'd10820};
                15'd12875 : data_rom <= {16'd30931, 16'd10817};
                15'd12876 : data_rom <= {16'd30932, 16'd10814};
                15'd12877 : data_rom <= {16'd30933, 16'd10811};
                15'd12878 : data_rom <= {16'd30934, 16'd10808};
                15'd12879 : data_rom <= {16'd30935, 16'd10805};
                15'd12880 : data_rom <= {16'd30936, 16'd10802};
                15'd12881 : data_rom <= {16'd30937, 16'd10799};
                15'd12882 : data_rom <= {16'd30938, 16'd10796};
                15'd12883 : data_rom <= {16'd30939, 16'd10793};
                15'd12884 : data_rom <= {16'd30940, 16'd10790};
                15'd12885 : data_rom <= {16'd30941, 16'd10787};
                15'd12886 : data_rom <= {16'd30942, 16'd10784};
                15'd12887 : data_rom <= {16'd30943, 16'd10781};
                15'd12888 : data_rom <= {16'd30944, 16'd10778};
                15'd12889 : data_rom <= {16'd30945, 16'd10775};
                15'd12890 : data_rom <= {16'd30946, 16'd10772};
                15'd12891 : data_rom <= {16'd30947, 16'd10769};
                15'd12892 : data_rom <= {16'd30948, 16'd10766};
                15'd12893 : data_rom <= {16'd30949, 16'd10763};
                15'd12894 : data_rom <= {16'd30950, 16'd10760};
                15'd12895 : data_rom <= {16'd30951, 16'd10757};
                15'd12896 : data_rom <= {16'd30952, 16'd10754};
                15'd12897 : data_rom <= {16'd30953, 16'd10751};
                15'd12898 : data_rom <= {16'd30954, 16'd10748};
                15'd12899 : data_rom <= {16'd30955, 16'd10745};
                15'd12900 : data_rom <= {16'd30956, 16'd10742};
                15'd12901 : data_rom <= {16'd30957, 16'd10739};
                15'd12902 : data_rom <= {16'd30958, 16'd10737};
                15'd12903 : data_rom <= {16'd30960, 16'd10734};
                15'd12904 : data_rom <= {16'd30961, 16'd10731};
                15'd12905 : data_rom <= {16'd30962, 16'd10728};
                15'd12906 : data_rom <= {16'd30963, 16'd10725};
                15'd12907 : data_rom <= {16'd30964, 16'd10722};
                15'd12908 : data_rom <= {16'd30965, 16'd10719};
                15'd12909 : data_rom <= {16'd30966, 16'd10716};
                15'd12910 : data_rom <= {16'd30967, 16'd10713};
                15'd12911 : data_rom <= {16'd30968, 16'd10710};
                15'd12912 : data_rom <= {16'd30969, 16'd10707};
                15'd12913 : data_rom <= {16'd30970, 16'd10704};
                15'd12914 : data_rom <= {16'd30971, 16'd10701};
                15'd12915 : data_rom <= {16'd30972, 16'd10698};
                15'd12916 : data_rom <= {16'd30973, 16'd10695};
                15'd12917 : data_rom <= {16'd30974, 16'd10692};
                15'd12918 : data_rom <= {16'd30975, 16'd10689};
                15'd12919 : data_rom <= {16'd30976, 16'd10686};
                15'd12920 : data_rom <= {16'd30977, 16'd10683};
                15'd12921 : data_rom <= {16'd30978, 16'd10680};
                15'd12922 : data_rom <= {16'd30979, 16'd10677};
                15'd12923 : data_rom <= {16'd30980, 16'd10674};
                15'd12924 : data_rom <= {16'd30981, 16'd10671};
                15'd12925 : data_rom <= {16'd30982, 16'd10668};
                15'd12926 : data_rom <= {16'd30983, 16'd10665};
                15'd12927 : data_rom <= {16'd30984, 16'd10662};
                15'd12928 : data_rom <= {16'd30985, 16'd10659};
                15'd12929 : data_rom <= {16'd30986, 16'd10656};
                15'd12930 : data_rom <= {16'd30987, 16'd10653};
                15'd12931 : data_rom <= {16'd30988, 16'd10650};
                15'd12932 : data_rom <= {16'd30989, 16'd10647};
                15'd12933 : data_rom <= {16'd30990, 16'd10644};
                15'd12934 : data_rom <= {16'd30991, 16'd10641};
                15'd12935 : data_rom <= {16'd30992, 16'd10639};
                15'd12936 : data_rom <= {16'd30993, 16'd10636};
                15'd12937 : data_rom <= {16'd30994, 16'd10633};
                15'd12938 : data_rom <= {16'd30995, 16'd10630};
                15'd12939 : data_rom <= {16'd30996, 16'd10627};
                15'd12940 : data_rom <= {16'd30997, 16'd10624};
                15'd12941 : data_rom <= {16'd30998, 16'd10621};
                15'd12942 : data_rom <= {16'd30999, 16'd10618};
                15'd12943 : data_rom <= {16'd31000, 16'd10615};
                15'd12944 : data_rom <= {16'd31001, 16'd10612};
                15'd12945 : data_rom <= {16'd31002, 16'd10609};
                15'd12946 : data_rom <= {16'd31003, 16'd10606};
                15'd12947 : data_rom <= {16'd31005, 16'd10603};
                15'd12948 : data_rom <= {16'd31006, 16'd10600};
                15'd12949 : data_rom <= {16'd31007, 16'd10597};
                15'd12950 : data_rom <= {16'd31008, 16'd10594};
                15'd12951 : data_rom <= {16'd31009, 16'd10591};
                15'd12952 : data_rom <= {16'd31010, 16'd10588};
                15'd12953 : data_rom <= {16'd31011, 16'd10585};
                15'd12954 : data_rom <= {16'd31012, 16'd10582};
                15'd12955 : data_rom <= {16'd31013, 16'd10579};
                15'd12956 : data_rom <= {16'd31014, 16'd10576};
                15'd12957 : data_rom <= {16'd31015, 16'd10573};
                15'd12958 : data_rom <= {16'd31016, 16'd10570};
                15'd12959 : data_rom <= {16'd31017, 16'd10567};
                15'd12960 : data_rom <= {16'd31018, 16'd10564};
                15'd12961 : data_rom <= {16'd31019, 16'd10561};
                15'd12962 : data_rom <= {16'd31020, 16'd10558};
                15'd12963 : data_rom <= {16'd31021, 16'd10555};
                15'd12964 : data_rom <= {16'd31022, 16'd10552};
                15'd12965 : data_rom <= {16'd31023, 16'd10549};
                15'd12966 : data_rom <= {16'd31024, 16'd10546};
                15'd12967 : data_rom <= {16'd31025, 16'd10543};
                15'd12968 : data_rom <= {16'd31026, 16'd10540};
                15'd12969 : data_rom <= {16'd31027, 16'd10537};
                15'd12970 : data_rom <= {16'd31028, 16'd10534};
                15'd12971 : data_rom <= {16'd31029, 16'd10531};
                15'd12972 : data_rom <= {16'd31030, 16'd10528};
                15'd12973 : data_rom <= {16'd31031, 16'd10526};
                15'd12974 : data_rom <= {16'd31032, 16'd10523};
                15'd12975 : data_rom <= {16'd31033, 16'd10520};
                15'd12976 : data_rom <= {16'd31034, 16'd10517};
                15'd12977 : data_rom <= {16'd31035, 16'd10514};
                15'd12978 : data_rom <= {16'd31036, 16'd10511};
                15'd12979 : data_rom <= {16'd31037, 16'd10508};
                15'd12980 : data_rom <= {16'd31038, 16'd10505};
                15'd12981 : data_rom <= {16'd31039, 16'd10502};
                15'd12982 : data_rom <= {16'd31040, 16'd10499};
                15'd12983 : data_rom <= {16'd31041, 16'd10496};
                15'd12984 : data_rom <= {16'd31042, 16'd10493};
                15'd12985 : data_rom <= {16'd31043, 16'd10490};
                15'd12986 : data_rom <= {16'd31044, 16'd10487};
                15'd12987 : data_rom <= {16'd31045, 16'd10484};
                15'd12988 : data_rom <= {16'd31046, 16'd10481};
                15'd12989 : data_rom <= {16'd31047, 16'd10478};
                15'd12990 : data_rom <= {16'd31048, 16'd10475};
                15'd12991 : data_rom <= {16'd31049, 16'd10472};
                15'd12992 : data_rom <= {16'd31050, 16'd10469};
                15'd12993 : data_rom <= {16'd31051, 16'd10466};
                15'd12994 : data_rom <= {16'd31052, 16'd10463};
                15'd12995 : data_rom <= {16'd31053, 16'd10460};
                15'd12996 : data_rom <= {16'd31054, 16'd10457};
                15'd12997 : data_rom <= {16'd31055, 16'd10454};
                15'd12998 : data_rom <= {16'd31056, 16'd10451};
                15'd12999 : data_rom <= {16'd31057, 16'd10448};
                15'd13000 : data_rom <= {16'd31058, 16'd10445};
                15'd13001 : data_rom <= {16'd31059, 16'd10442};
                15'd13002 : data_rom <= {16'd31060, 16'd10439};
                15'd13003 : data_rom <= {16'd31061, 16'd10436};
                15'd13004 : data_rom <= {16'd31062, 16'd10433};
                15'd13005 : data_rom <= {16'd31063, 16'd10430};
                15'd13006 : data_rom <= {16'd31064, 16'd10427};
                15'd13007 : data_rom <= {16'd31065, 16'd10424};
                15'd13008 : data_rom <= {16'd31066, 16'd10421};
                15'd13009 : data_rom <= {16'd31067, 16'd10418};
                15'd13010 : data_rom <= {16'd31068, 16'd10415};
                15'd13011 : data_rom <= {16'd31069, 16'd10412};
                15'd13012 : data_rom <= {16'd31070, 16'd10409};
                15'd13013 : data_rom <= {16'd31071, 16'd10406};
                15'd13014 : data_rom <= {16'd31072, 16'd10403};
                15'd13015 : data_rom <= {16'd31073, 16'd10400};
                15'd13016 : data_rom <= {16'd31074, 16'd10398};
                15'd13017 : data_rom <= {16'd31075, 16'd10395};
                15'd13018 : data_rom <= {16'd31076, 16'd10392};
                15'd13019 : data_rom <= {16'd31077, 16'd10389};
                15'd13020 : data_rom <= {16'd31078, 16'd10386};
                15'd13021 : data_rom <= {16'd31079, 16'd10383};
                15'd13022 : data_rom <= {16'd31080, 16'd10380};
                15'd13023 : data_rom <= {16'd31081, 16'd10377};
                15'd13024 : data_rom <= {16'd31082, 16'd10374};
                15'd13025 : data_rom <= {16'd31083, 16'd10371};
                15'd13026 : data_rom <= {16'd31084, 16'd10368};
                15'd13027 : data_rom <= {16'd31085, 16'd10365};
                15'd13028 : data_rom <= {16'd31086, 16'd10362};
                15'd13029 : data_rom <= {16'd31087, 16'd10359};
                15'd13030 : data_rom <= {16'd31088, 16'd10356};
                15'd13031 : data_rom <= {16'd31089, 16'd10353};
                15'd13032 : data_rom <= {16'd31090, 16'd10350};
                15'd13033 : data_rom <= {16'd31091, 16'd10347};
                15'd13034 : data_rom <= {16'd31092, 16'd10344};
                15'd13035 : data_rom <= {16'd31093, 16'd10341};
                15'd13036 : data_rom <= {16'd31094, 16'd10338};
                15'd13037 : data_rom <= {16'd31095, 16'd10335};
                15'd13038 : data_rom <= {16'd31096, 16'd10332};
                15'd13039 : data_rom <= {16'd31097, 16'd10329};
                15'd13040 : data_rom <= {16'd31098, 16'd10326};
                15'd13041 : data_rom <= {16'd31099, 16'd10323};
                15'd13042 : data_rom <= {16'd31100, 16'd10320};
                15'd13043 : data_rom <= {16'd31101, 16'd10317};
                15'd13044 : data_rom <= {16'd31102, 16'd10314};
                15'd13045 : data_rom <= {16'd31103, 16'd10311};
                15'd13046 : data_rom <= {16'd31104, 16'd10308};
                15'd13047 : data_rom <= {16'd31105, 16'd10305};
                15'd13048 : data_rom <= {16'd31106, 16'd10302};
                15'd13049 : data_rom <= {16'd31107, 16'd10299};
                15'd13050 : data_rom <= {16'd31108, 16'd10296};
                15'd13051 : data_rom <= {16'd31109, 16'd10293};
                15'd13052 : data_rom <= {16'd31110, 16'd10290};
                15'd13053 : data_rom <= {16'd31111, 16'd10287};
                15'd13054 : data_rom <= {16'd31112, 16'd10284};
                15'd13055 : data_rom <= {16'd31113, 16'd10281};
                15'd13056 : data_rom <= {16'd31114, 16'd10278};
                15'd13057 : data_rom <= {16'd31115, 16'd10275};
                15'd13058 : data_rom <= {16'd31116, 16'd10272};
                15'd13059 : data_rom <= {16'd31117, 16'd10269};
                15'd13060 : data_rom <= {16'd31118, 16'd10266};
                15'd13061 : data_rom <= {16'd31119, 16'd10263};
                15'd13062 : data_rom <= {16'd31120, 16'd10260};
                15'd13063 : data_rom <= {16'd31121, 16'd10257};
                15'd13064 : data_rom <= {16'd31122, 16'd10254};
                15'd13065 : data_rom <= {16'd31122, 16'd10251};
                15'd13066 : data_rom <= {16'd31123, 16'd10248};
                15'd13067 : data_rom <= {16'd31124, 16'd10245};
                15'd13068 : data_rom <= {16'd31125, 16'd10242};
                15'd13069 : data_rom <= {16'd31126, 16'd10239};
                15'd13070 : data_rom <= {16'd31127, 16'd10236};
                15'd13071 : data_rom <= {16'd31128, 16'd10234};
                15'd13072 : data_rom <= {16'd31129, 16'd10231};
                15'd13073 : data_rom <= {16'd31130, 16'd10228};
                15'd13074 : data_rom <= {16'd31131, 16'd10225};
                15'd13075 : data_rom <= {16'd31132, 16'd10222};
                15'd13076 : data_rom <= {16'd31133, 16'd10219};
                15'd13077 : data_rom <= {16'd31134, 16'd10216};
                15'd13078 : data_rom <= {16'd31135, 16'd10213};
                15'd13079 : data_rom <= {16'd31136, 16'd10210};
                15'd13080 : data_rom <= {16'd31137, 16'd10207};
                15'd13081 : data_rom <= {16'd31138, 16'd10204};
                15'd13082 : data_rom <= {16'd31139, 16'd10201};
                15'd13083 : data_rom <= {16'd31140, 16'd10198};
                15'd13084 : data_rom <= {16'd31141, 16'd10195};
                15'd13085 : data_rom <= {16'd31142, 16'd10192};
                15'd13086 : data_rom <= {16'd31143, 16'd10189};
                15'd13087 : data_rom <= {16'd31144, 16'd10186};
                15'd13088 : data_rom <= {16'd31145, 16'd10183};
                15'd13089 : data_rom <= {16'd31146, 16'd10180};
                15'd13090 : data_rom <= {16'd31147, 16'd10177};
                15'd13091 : data_rom <= {16'd31148, 16'd10174};
                15'd13092 : data_rom <= {16'd31149, 16'd10171};
                15'd13093 : data_rom <= {16'd31150, 16'd10168};
                15'd13094 : data_rom <= {16'd31151, 16'd10165};
                15'd13095 : data_rom <= {16'd31152, 16'd10162};
                15'd13096 : data_rom <= {16'd31153, 16'd10159};
                15'd13097 : data_rom <= {16'd31154, 16'd10156};
                15'd13098 : data_rom <= {16'd31155, 16'd10153};
                15'd13099 : data_rom <= {16'd31156, 16'd10150};
                15'd13100 : data_rom <= {16'd31157, 16'd10147};
                15'd13101 : data_rom <= {16'd31158, 16'd10144};
                15'd13102 : data_rom <= {16'd31159, 16'd10141};
                15'd13103 : data_rom <= {16'd31160, 16'd10138};
                15'd13104 : data_rom <= {16'd31161, 16'd10135};
                15'd13105 : data_rom <= {16'd31162, 16'd10132};
                15'd13106 : data_rom <= {16'd31163, 16'd10129};
                15'd13107 : data_rom <= {16'd31164, 16'd10126};
                15'd13108 : data_rom <= {16'd31164, 16'd10123};
                15'd13109 : data_rom <= {16'd31165, 16'd10120};
                15'd13110 : data_rom <= {16'd31166, 16'd10117};
                15'd13111 : data_rom <= {16'd31167, 16'd10114};
                15'd13112 : data_rom <= {16'd31168, 16'd10111};
                15'd13113 : data_rom <= {16'd31169, 16'd10108};
                15'd13114 : data_rom <= {16'd31170, 16'd10105};
                15'd13115 : data_rom <= {16'd31171, 16'd10102};
                15'd13116 : data_rom <= {16'd31172, 16'd10099};
                15'd13117 : data_rom <= {16'd31173, 16'd10096};
                15'd13118 : data_rom <= {16'd31174, 16'd10093};
                15'd13119 : data_rom <= {16'd31175, 16'd10090};
                15'd13120 : data_rom <= {16'd31176, 16'd10087};
                15'd13121 : data_rom <= {16'd31177, 16'd10084};
                15'd13122 : data_rom <= {16'd31178, 16'd10081};
                15'd13123 : data_rom <= {16'd31179, 16'd10078};
                15'd13124 : data_rom <= {16'd31180, 16'd10075};
                15'd13125 : data_rom <= {16'd31181, 16'd10072};
                15'd13126 : data_rom <= {16'd31182, 16'd10069};
                15'd13127 : data_rom <= {16'd31183, 16'd10066};
                15'd13128 : data_rom <= {16'd31184, 16'd10063};
                15'd13129 : data_rom <= {16'd31185, 16'd10060};
                15'd13130 : data_rom <= {16'd31186, 16'd10057};
                15'd13131 : data_rom <= {16'd31187, 16'd10054};
                15'd13132 : data_rom <= {16'd31188, 16'd10051};
                15'd13133 : data_rom <= {16'd31189, 16'd10048};
                15'd13134 : data_rom <= {16'd31190, 16'd10045};
                15'd13135 : data_rom <= {16'd31191, 16'd10042};
                15'd13136 : data_rom <= {16'd31192, 16'd10039};
                15'd13137 : data_rom <= {16'd31193, 16'd10036};
                15'd13138 : data_rom <= {16'd31193, 16'd10033};
                15'd13139 : data_rom <= {16'd31194, 16'd10030};
                15'd13140 : data_rom <= {16'd31195, 16'd10027};
                15'd13141 : data_rom <= {16'd31196, 16'd10024};
                15'd13142 : data_rom <= {16'd31197, 16'd10021};
                15'd13143 : data_rom <= {16'd31198, 16'd10018};
                15'd13144 : data_rom <= {16'd31199, 16'd10015};
                15'd13145 : data_rom <= {16'd31200, 16'd10012};
                15'd13146 : data_rom <= {16'd31201, 16'd10009};
                15'd13147 : data_rom <= {16'd31202, 16'd10006};
                15'd13148 : data_rom <= {16'd31203, 16'd10003};
                15'd13149 : data_rom <= {16'd31204, 16'd10000};
                15'd13150 : data_rom <= {16'd31205, 16'd9997};
                15'd13151 : data_rom <= {16'd31206, 16'd9994};
                15'd13152 : data_rom <= {16'd31207, 16'd9991};
                15'd13153 : data_rom <= {16'd31208, 16'd9988};
                15'd13154 : data_rom <= {16'd31209, 16'd9985};
                15'd13155 : data_rom <= {16'd31210, 16'd9982};
                15'd13156 : data_rom <= {16'd31211, 16'd9979};
                15'd13157 : data_rom <= {16'd31212, 16'd9976};
                15'd13158 : data_rom <= {16'd31213, 16'd9974};
                15'd13159 : data_rom <= {16'd31214, 16'd9971};
                15'd13160 : data_rom <= {16'd31215, 16'd9968};
                15'd13161 : data_rom <= {16'd31216, 16'd9965};
                15'd13162 : data_rom <= {16'd31216, 16'd9962};
                15'd13163 : data_rom <= {16'd31217, 16'd9959};
                15'd13164 : data_rom <= {16'd31218, 16'd9956};
                15'd13165 : data_rom <= {16'd31219, 16'd9953};
                15'd13166 : data_rom <= {16'd31220, 16'd9950};
                15'd13167 : data_rom <= {16'd31221, 16'd9947};
                15'd13168 : data_rom <= {16'd31222, 16'd9944};
                15'd13169 : data_rom <= {16'd31223, 16'd9941};
                15'd13170 : data_rom <= {16'd31224, 16'd9938};
                15'd13171 : data_rom <= {16'd31225, 16'd9935};
                15'd13172 : data_rom <= {16'd31226, 16'd9932};
                15'd13173 : data_rom <= {16'd31227, 16'd9929};
                15'd13174 : data_rom <= {16'd31228, 16'd9926};
                15'd13175 : data_rom <= {16'd31229, 16'd9923};
                15'd13176 : data_rom <= {16'd31230, 16'd9920};
                15'd13177 : data_rom <= {16'd31231, 16'd9917};
                15'd13178 : data_rom <= {16'd31232, 16'd9914};
                15'd13179 : data_rom <= {16'd31233, 16'd9911};
                15'd13180 : data_rom <= {16'd31234, 16'd9908};
                15'd13181 : data_rom <= {16'd31235, 16'd9905};
                15'd13182 : data_rom <= {16'd31236, 16'd9902};
                15'd13183 : data_rom <= {16'd31236, 16'd9899};
                15'd13184 : data_rom <= {16'd31237, 16'd9896};
                15'd13185 : data_rom <= {16'd31238, 16'd9893};
                15'd13186 : data_rom <= {16'd31239, 16'd9890};
                15'd13187 : data_rom <= {16'd31240, 16'd9887};
                15'd13188 : data_rom <= {16'd31241, 16'd9884};
                15'd13189 : data_rom <= {16'd31242, 16'd9881};
                15'd13190 : data_rom <= {16'd31243, 16'd9878};
                15'd13191 : data_rom <= {16'd31244, 16'd9875};
                15'd13192 : data_rom <= {16'd31245, 16'd9872};
                15'd13193 : data_rom <= {16'd31246, 16'd9869};
                15'd13194 : data_rom <= {16'd31247, 16'd9866};
                15'd13195 : data_rom <= {16'd31248, 16'd9863};
                15'd13196 : data_rom <= {16'd31249, 16'd9860};
                15'd13197 : data_rom <= {16'd31250, 16'd9857};
                15'd13198 : data_rom <= {16'd31251, 16'd9854};
                15'd13199 : data_rom <= {16'd31252, 16'd9851};
                15'd13200 : data_rom <= {16'd31253, 16'd9848};
                15'd13201 : data_rom <= {16'd31254, 16'd9845};
                15'd13202 : data_rom <= {16'd31254, 16'd9842};
                15'd13203 : data_rom <= {16'd31255, 16'd9839};
                15'd13204 : data_rom <= {16'd31256, 16'd9836};
                15'd13205 : data_rom <= {16'd31257, 16'd9833};
                15'd13206 : data_rom <= {16'd31258, 16'd9830};
                15'd13207 : data_rom <= {16'd31259, 16'd9827};
                15'd13208 : data_rom <= {16'd31260, 16'd9824};
                15'd13209 : data_rom <= {16'd31261, 16'd9821};
                15'd13210 : data_rom <= {16'd31262, 16'd9818};
                15'd13211 : data_rom <= {16'd31263, 16'd9815};
                15'd13212 : data_rom <= {16'd31264, 16'd9812};
                15'd13213 : data_rom <= {16'd31265, 16'd9809};
                15'd13214 : data_rom <= {16'd31266, 16'd9806};
                15'd13215 : data_rom <= {16'd31267, 16'd9803};
                15'd13216 : data_rom <= {16'd31268, 16'd9800};
                15'd13217 : data_rom <= {16'd31269, 16'd9797};
                15'd13218 : data_rom <= {16'd31270, 16'd9794};
                15'd13219 : data_rom <= {16'd31270, 16'd9791};
                15'd13220 : data_rom <= {16'd31271, 16'd9788};
                15'd13221 : data_rom <= {16'd31272, 16'd9785};
                15'd13222 : data_rom <= {16'd31273, 16'd9782};
                15'd13223 : data_rom <= {16'd31274, 16'd9779};
                15'd13224 : data_rom <= {16'd31275, 16'd9776};
                15'd13225 : data_rom <= {16'd31276, 16'd9773};
                15'd13226 : data_rom <= {16'd31277, 16'd9770};
                15'd13227 : data_rom <= {16'd31278, 16'd9767};
                15'd13228 : data_rom <= {16'd31279, 16'd9764};
                15'd13229 : data_rom <= {16'd31280, 16'd9761};
                15'd13230 : data_rom <= {16'd31281, 16'd9758};
                15'd13231 : data_rom <= {16'd31282, 16'd9755};
                15'd13232 : data_rom <= {16'd31283, 16'd9752};
                15'd13233 : data_rom <= {16'd31284, 16'd9749};
                15'd13234 : data_rom <= {16'd31285, 16'd9746};
                15'd13235 : data_rom <= {16'd31285, 16'd9743};
                15'd13236 : data_rom <= {16'd31286, 16'd9740};
                15'd13237 : data_rom <= {16'd31287, 16'd9737};
                15'd13238 : data_rom <= {16'd31288, 16'd9734};
                15'd13239 : data_rom <= {16'd31289, 16'd9731};
                15'd13240 : data_rom <= {16'd31290, 16'd9728};
                15'd13241 : data_rom <= {16'd31291, 16'd9725};
                15'd13242 : data_rom <= {16'd31292, 16'd9722};
                15'd13243 : data_rom <= {16'd31293, 16'd9719};
                15'd13244 : data_rom <= {16'd31294, 16'd9716};
                15'd13245 : data_rom <= {16'd31295, 16'd9713};
                15'd13246 : data_rom <= {16'd31296, 16'd9710};
                15'd13247 : data_rom <= {16'd31297, 16'd9707};
                15'd13248 : data_rom <= {16'd31298, 16'd9704};
                15'd13249 : data_rom <= {16'd31298, 16'd9701};
                15'd13250 : data_rom <= {16'd31299, 16'd9698};
                15'd13251 : data_rom <= {16'd31300, 16'd9695};
                15'd13252 : data_rom <= {16'd31301, 16'd9692};
                15'd13253 : data_rom <= {16'd31302, 16'd9689};
                15'd13254 : data_rom <= {16'd31303, 16'd9686};
                15'd13255 : data_rom <= {16'd31304, 16'd9683};
                15'd13256 : data_rom <= {16'd31305, 16'd9680};
                15'd13257 : data_rom <= {16'd31306, 16'd9677};
                15'd13258 : data_rom <= {16'd31307, 16'd9674};
                15'd13259 : data_rom <= {16'd31308, 16'd9671};
                15'd13260 : data_rom <= {16'd31309, 16'd9668};
                15'd13261 : data_rom <= {16'd31310, 16'd9665};
                15'd13262 : data_rom <= {16'd31311, 16'd9662};
                15'd13263 : data_rom <= {16'd31311, 16'd9659};
                15'd13264 : data_rom <= {16'd31312, 16'd9656};
                15'd13265 : data_rom <= {16'd31313, 16'd9653};
                15'd13266 : data_rom <= {16'd31314, 16'd9650};
                15'd13267 : data_rom <= {16'd31315, 16'd9647};
                15'd13268 : data_rom <= {16'd31316, 16'd9644};
                15'd13269 : data_rom <= {16'd31317, 16'd9641};
                15'd13270 : data_rom <= {16'd31318, 16'd9638};
                15'd13271 : data_rom <= {16'd31319, 16'd9635};
                15'd13272 : data_rom <= {16'd31320, 16'd9632};
                15'd13273 : data_rom <= {16'd31321, 16'd9629};
                15'd13274 : data_rom <= {16'd31322, 16'd9626};
                15'd13275 : data_rom <= {16'd31323, 16'd9623};
                15'd13276 : data_rom <= {16'd31323, 16'd9620};
                15'd13277 : data_rom <= {16'd31324, 16'd9617};
                15'd13278 : data_rom <= {16'd31325, 16'd9614};
                15'd13279 : data_rom <= {16'd31326, 16'd9611};
                15'd13280 : data_rom <= {16'd31327, 16'd9608};
                15'd13281 : data_rom <= {16'd31328, 16'd9605};
                15'd13282 : data_rom <= {16'd31329, 16'd9602};
                15'd13283 : data_rom <= {16'd31330, 16'd9599};
                15'd13284 : data_rom <= {16'd31331, 16'd9596};
                15'd13285 : data_rom <= {16'd31332, 16'd9593};
                15'd13286 : data_rom <= {16'd31333, 16'd9590};
                15'd13287 : data_rom <= {16'd31334, 16'd9587};
                15'd13288 : data_rom <= {16'd31335, 16'd9584};
                15'd13289 : data_rom <= {16'd31335, 16'd9581};
                15'd13290 : data_rom <= {16'd31336, 16'd9578};
                15'd13291 : data_rom <= {16'd31337, 16'd9575};
                15'd13292 : data_rom <= {16'd31338, 16'd9572};
                15'd13293 : data_rom <= {16'd31339, 16'd9569};
                15'd13294 : data_rom <= {16'd31340, 16'd9566};
                15'd13295 : data_rom <= {16'd31341, 16'd9563};
                15'd13296 : data_rom <= {16'd31342, 16'd9560};
                15'd13297 : data_rom <= {16'd31343, 16'd9557};
                15'd13298 : data_rom <= {16'd31344, 16'd9554};
                15'd13299 : data_rom <= {16'd31345, 16'd9551};
                15'd13300 : data_rom <= {16'd31346, 16'd9548};
                15'd13301 : data_rom <= {16'd31346, 16'd9545};
                15'd13302 : data_rom <= {16'd31347, 16'd9542};
                15'd13303 : data_rom <= {16'd31348, 16'd9539};
                15'd13304 : data_rom <= {16'd31349, 16'd9536};
                15'd13305 : data_rom <= {16'd31350, 16'd9533};
                15'd13306 : data_rom <= {16'd31351, 16'd9530};
                15'd13307 : data_rom <= {16'd31352, 16'd9527};
                15'd13308 : data_rom <= {16'd31353, 16'd9524};
                15'd13309 : data_rom <= {16'd31354, 16'd9521};
                15'd13310 : data_rom <= {16'd31355, 16'd9518};
                15'd13311 : data_rom <= {16'd31356, 16'd9515};
                15'd13312 : data_rom <= {16'd31357, 16'd9512};
                15'd13313 : data_rom <= {16'd31357, 16'd9509};
                15'd13314 : data_rom <= {16'd31358, 16'd9506};
                15'd13315 : data_rom <= {16'd31359, 16'd9503};
                15'd13316 : data_rom <= {16'd31360, 16'd9500};
                15'd13317 : data_rom <= {16'd31361, 16'd9497};
                15'd13318 : data_rom <= {16'd31362, 16'd9494};
                15'd13319 : data_rom <= {16'd31363, 16'd9491};
                15'd13320 : data_rom <= {16'd31364, 16'd9488};
                15'd13321 : data_rom <= {16'd31365, 16'd9485};
                15'd13322 : data_rom <= {16'd31366, 16'd9482};
                15'd13323 : data_rom <= {16'd31367, 16'd9479};
                15'd13324 : data_rom <= {16'd31367, 16'd9476};
                15'd13325 : data_rom <= {16'd31368, 16'd9472};
                15'd13326 : data_rom <= {16'd31369, 16'd9469};
                15'd13327 : data_rom <= {16'd31370, 16'd9466};
                15'd13328 : data_rom <= {16'd31371, 16'd9463};
                15'd13329 : data_rom <= {16'd31372, 16'd9460};
                15'd13330 : data_rom <= {16'd31373, 16'd9457};
                15'd13331 : data_rom <= {16'd31374, 16'd9454};
                15'd13332 : data_rom <= {16'd31375, 16'd9451};
                15'd13333 : data_rom <= {16'd31376, 16'd9448};
                15'd13334 : data_rom <= {16'd31377, 16'd9445};
                15'd13335 : data_rom <= {16'd31377, 16'd9442};
                15'd13336 : data_rom <= {16'd31378, 16'd9439};
                15'd13337 : data_rom <= {16'd31379, 16'd9436};
                15'd13338 : data_rom <= {16'd31380, 16'd9433};
                15'd13339 : data_rom <= {16'd31381, 16'd9430};
                15'd13340 : data_rom <= {16'd31382, 16'd9427};
                15'd13341 : data_rom <= {16'd31383, 16'd9424};
                15'd13342 : data_rom <= {16'd31384, 16'd9421};
                15'd13343 : data_rom <= {16'd31385, 16'd9418};
                15'd13344 : data_rom <= {16'd31386, 16'd9415};
                15'd13345 : data_rom <= {16'd31386, 16'd9412};
                15'd13346 : data_rom <= {16'd31387, 16'd9409};
                15'd13347 : data_rom <= {16'd31388, 16'd9406};
                15'd13348 : data_rom <= {16'd31389, 16'd9403};
                15'd13349 : data_rom <= {16'd31390, 16'd9400};
                15'd13350 : data_rom <= {16'd31391, 16'd9397};
                15'd13351 : data_rom <= {16'd31392, 16'd9394};
                15'd13352 : data_rom <= {16'd31393, 16'd9391};
                15'd13353 : data_rom <= {16'd31394, 16'd9388};
                15'd13354 : data_rom <= {16'd31395, 16'd9385};
                15'd13355 : data_rom <= {16'd31395, 16'd9382};
                15'd13356 : data_rom <= {16'd31396, 16'd9379};
                15'd13357 : data_rom <= {16'd31397, 16'd9376};
                15'd13358 : data_rom <= {16'd31398, 16'd9373};
                15'd13359 : data_rom <= {16'd31399, 16'd9370};
                15'd13360 : data_rom <= {16'd31400, 16'd9367};
                15'd13361 : data_rom <= {16'd31401, 16'd9364};
                15'd13362 : data_rom <= {16'd31402, 16'd9361};
                15'd13363 : data_rom <= {16'd31403, 16'd9358};
                15'd13364 : data_rom <= {16'd31404, 16'd9355};
                15'd13365 : data_rom <= {16'd31404, 16'd9352};
                15'd13366 : data_rom <= {16'd31405, 16'd9349};
                15'd13367 : data_rom <= {16'd31406, 16'd9346};
                15'd13368 : data_rom <= {16'd31407, 16'd9343};
                15'd13369 : data_rom <= {16'd31408, 16'd9340};
                15'd13370 : data_rom <= {16'd31409, 16'd9337};
                15'd13371 : data_rom <= {16'd31410, 16'd9334};
                15'd13372 : data_rom <= {16'd31411, 16'd9331};
                15'd13373 : data_rom <= {16'd31412, 16'd9328};
                15'd13374 : data_rom <= {16'd31412, 16'd9325};
                15'd13375 : data_rom <= {16'd31413, 16'd9322};
                15'd13376 : data_rom <= {16'd31414, 16'd9319};
                15'd13377 : data_rom <= {16'd31415, 16'd9316};
                15'd13378 : data_rom <= {16'd31416, 16'd9313};
                15'd13379 : data_rom <= {16'd31417, 16'd9310};
                15'd13380 : data_rom <= {16'd31418, 16'd9307};
                15'd13381 : data_rom <= {16'd31419, 16'd9304};
                15'd13382 : data_rom <= {16'd31420, 16'd9301};
                15'd13383 : data_rom <= {16'd31421, 16'd9298};
                15'd13384 : data_rom <= {16'd31421, 16'd9295};
                15'd13385 : data_rom <= {16'd31422, 16'd9292};
                15'd13386 : data_rom <= {16'd31423, 16'd9289};
                15'd13387 : data_rom <= {16'd31424, 16'd9286};
                15'd13388 : data_rom <= {16'd31425, 16'd9283};
                15'd13389 : data_rom <= {16'd31426, 16'd9280};
                15'd13390 : data_rom <= {16'd31427, 16'd9277};
                15'd13391 : data_rom <= {16'd31428, 16'd9274};
                15'd13392 : data_rom <= {16'd31429, 16'd9271};
                15'd13393 : data_rom <= {16'd31429, 16'd9268};
                15'd13394 : data_rom <= {16'd31430, 16'd9265};
                15'd13395 : data_rom <= {16'd31431, 16'd9262};
                15'd13396 : data_rom <= {16'd31432, 16'd9259};
                15'd13397 : data_rom <= {16'd31433, 16'd9256};
                15'd13398 : data_rom <= {16'd31434, 16'd9253};
                15'd13399 : data_rom <= {16'd31435, 16'd9250};
                15'd13400 : data_rom <= {16'd31436, 16'd9247};
                15'd13401 : data_rom <= {16'd31437, 16'd9244};
                15'd13402 : data_rom <= {16'd31437, 16'd9241};
                15'd13403 : data_rom <= {16'd31438, 16'd9238};
                15'd13404 : data_rom <= {16'd31439, 16'd9235};
                15'd13405 : data_rom <= {16'd31440, 16'd9232};
                15'd13406 : data_rom <= {16'd31441, 16'd9229};
                15'd13407 : data_rom <= {16'd31442, 16'd9226};
                15'd13408 : data_rom <= {16'd31443, 16'd9223};
                15'd13409 : data_rom <= {16'd31444, 16'd9220};
                15'd13410 : data_rom <= {16'd31444, 16'd9217};
                15'd13411 : data_rom <= {16'd31445, 16'd9214};
                15'd13412 : data_rom <= {16'd31446, 16'd9211};
                15'd13413 : data_rom <= {16'd31447, 16'd9208};
                15'd13414 : data_rom <= {16'd31448, 16'd9204};
                15'd13415 : data_rom <= {16'd31449, 16'd9201};
                15'd13416 : data_rom <= {16'd31450, 16'd9198};
                15'd13417 : data_rom <= {16'd31451, 16'd9195};
                15'd13418 : data_rom <= {16'd31452, 16'd9192};
                15'd13419 : data_rom <= {16'd31452, 16'd9189};
                15'd13420 : data_rom <= {16'd31453, 16'd9186};
                15'd13421 : data_rom <= {16'd31454, 16'd9183};
                15'd13422 : data_rom <= {16'd31455, 16'd9180};
                15'd13423 : data_rom <= {16'd31456, 16'd9177};
                15'd13424 : data_rom <= {16'd31457, 16'd9174};
                15'd13425 : data_rom <= {16'd31458, 16'd9171};
                15'd13426 : data_rom <= {16'd31459, 16'd9168};
                15'd13427 : data_rom <= {16'd31459, 16'd9165};
                15'd13428 : data_rom <= {16'd31460, 16'd9162};
                15'd13429 : data_rom <= {16'd31461, 16'd9159};
                15'd13430 : data_rom <= {16'd31462, 16'd9156};
                15'd13431 : data_rom <= {16'd31463, 16'd9153};
                15'd13432 : data_rom <= {16'd31464, 16'd9150};
                15'd13433 : data_rom <= {16'd31465, 16'd9147};
                15'd13434 : data_rom <= {16'd31466, 16'd9144};
                15'd13435 : data_rom <= {16'd31466, 16'd9141};
                15'd13436 : data_rom <= {16'd31467, 16'd9138};
                15'd13437 : data_rom <= {16'd31468, 16'd9135};
                15'd13438 : data_rom <= {16'd31469, 16'd9132};
                15'd13439 : data_rom <= {16'd31470, 16'd9129};
                15'd13440 : data_rom <= {16'd31471, 16'd9126};
                15'd13441 : data_rom <= {16'd31472, 16'd9123};
                15'd13442 : data_rom <= {16'd31473, 16'd9120};
                15'd13443 : data_rom <= {16'd31473, 16'd9117};
                15'd13444 : data_rom <= {16'd31474, 16'd9114};
                15'd13445 : data_rom <= {16'd31475, 16'd9111};
                15'd13446 : data_rom <= {16'd31476, 16'd9108};
                15'd13447 : data_rom <= {16'd31477, 16'd9105};
                15'd13448 : data_rom <= {16'd31478, 16'd9102};
                15'd13449 : data_rom <= {16'd31479, 16'd9099};
                15'd13450 : data_rom <= {16'd31480, 16'd9096};
                15'd13451 : data_rom <= {16'd31480, 16'd9093};
                15'd13452 : data_rom <= {16'd31481, 16'd9090};
                15'd13453 : data_rom <= {16'd31482, 16'd9087};
                15'd13454 : data_rom <= {16'd31483, 16'd9084};
                15'd13455 : data_rom <= {16'd31484, 16'd9081};
                15'd13456 : data_rom <= {16'd31485, 16'd9078};
                15'd13457 : data_rom <= {16'd31486, 16'd9075};
                15'd13458 : data_rom <= {16'd31487, 16'd9072};
                15'd13459 : data_rom <= {16'd31487, 16'd9069};
                15'd13460 : data_rom <= {16'd31488, 16'd9066};
                15'd13461 : data_rom <= {16'd31489, 16'd9063};
                15'd13462 : data_rom <= {16'd31490, 16'd9060};
                15'd13463 : data_rom <= {16'd31491, 16'd9057};
                15'd13464 : data_rom <= {16'd31492, 16'd9054};
                15'd13465 : data_rom <= {16'd31493, 16'd9051};
                15'd13466 : data_rom <= {16'd31494, 16'd9048};
                15'd13467 : data_rom <= {16'd31494, 16'd9045};
                15'd13468 : data_rom <= {16'd31495, 16'd9042};
                15'd13469 : data_rom <= {16'd31496, 16'd9039};
                15'd13470 : data_rom <= {16'd31497, 16'd9036};
                15'd13471 : data_rom <= {16'd31498, 16'd9032};
                15'd13472 : data_rom <= {16'd31499, 16'd9029};
                15'd13473 : data_rom <= {16'd31500, 16'd9026};
                15'd13474 : data_rom <= {16'd31500, 16'd9023};
                15'd13475 : data_rom <= {16'd31501, 16'd9020};
                15'd13476 : data_rom <= {16'd31502, 16'd9017};
                15'd13477 : data_rom <= {16'd31503, 16'd9014};
                15'd13478 : data_rom <= {16'd31504, 16'd9011};
                15'd13479 : data_rom <= {16'd31505, 16'd9008};
                15'd13480 : data_rom <= {16'd31506, 16'd9005};
                15'd13481 : data_rom <= {16'd31507, 16'd9002};
                15'd13482 : data_rom <= {16'd31507, 16'd8999};
                15'd13483 : data_rom <= {16'd31508, 16'd8996};
                15'd13484 : data_rom <= {16'd31509, 16'd8993};
                15'd13485 : data_rom <= {16'd31510, 16'd8990};
                15'd13486 : data_rom <= {16'd31511, 16'd8987};
                15'd13487 : data_rom <= {16'd31512, 16'd8984};
                15'd13488 : data_rom <= {16'd31513, 16'd8981};
                15'd13489 : data_rom <= {16'd31513, 16'd8978};
                15'd13490 : data_rom <= {16'd31514, 16'd8975};
                15'd13491 : data_rom <= {16'd31515, 16'd8972};
                15'd13492 : data_rom <= {16'd31516, 16'd8969};
                15'd13493 : data_rom <= {16'd31517, 16'd8966};
                15'd13494 : data_rom <= {16'd31518, 16'd8963};
                15'd13495 : data_rom <= {16'd31519, 16'd8960};
                15'd13496 : data_rom <= {16'd31519, 16'd8957};
                15'd13497 : data_rom <= {16'd31520, 16'd8954};
                15'd13498 : data_rom <= {16'd31521, 16'd8951};
                15'd13499 : data_rom <= {16'd31522, 16'd8948};
                15'd13500 : data_rom <= {16'd31523, 16'd8945};
                15'd13501 : data_rom <= {16'd31524, 16'd8942};
                15'd13502 : data_rom <= {16'd31525, 16'd8939};
                15'd13503 : data_rom <= {16'd31525, 16'd8936};
                15'd13504 : data_rom <= {16'd31526, 16'd8933};
                15'd13505 : data_rom <= {16'd31527, 16'd8930};
                15'd13506 : data_rom <= {16'd31528, 16'd8927};
                15'd13507 : data_rom <= {16'd31529, 16'd8924};
                15'd13508 : data_rom <= {16'd31530, 16'd8921};
                15'd13509 : data_rom <= {16'd31531, 16'd8918};
                15'd13510 : data_rom <= {16'd31531, 16'd8915};
                15'd13511 : data_rom <= {16'd31532, 16'd8912};
                15'd13512 : data_rom <= {16'd31533, 16'd8909};
                15'd13513 : data_rom <= {16'd31534, 16'd8906};
                15'd13514 : data_rom <= {16'd31535, 16'd8903};
                15'd13515 : data_rom <= {16'd31536, 16'd8900};
                15'd13516 : data_rom <= {16'd31537, 16'd8897};
                15'd13517 : data_rom <= {16'd31537, 16'd8893};
                15'd13518 : data_rom <= {16'd31538, 16'd8890};
                15'd13519 : data_rom <= {16'd31539, 16'd8887};
                15'd13520 : data_rom <= {16'd31540, 16'd8884};
                15'd13521 : data_rom <= {16'd31541, 16'd8881};
                15'd13522 : data_rom <= {16'd31542, 16'd8878};
                15'd13523 : data_rom <= {16'd31543, 16'd8875};
                15'd13524 : data_rom <= {16'd31543, 16'd8872};
                15'd13525 : data_rom <= {16'd31544, 16'd8869};
                15'd13526 : data_rom <= {16'd31545, 16'd8866};
                15'd13527 : data_rom <= {16'd31546, 16'd8863};
                15'd13528 : data_rom <= {16'd31547, 16'd8860};
                15'd13529 : data_rom <= {16'd31548, 16'd8857};
                15'd13530 : data_rom <= {16'd31548, 16'd8854};
                15'd13531 : data_rom <= {16'd31549, 16'd8851};
                15'd13532 : data_rom <= {16'd31550, 16'd8848};
                15'd13533 : data_rom <= {16'd31551, 16'd8845};
                15'd13534 : data_rom <= {16'd31552, 16'd8842};
                15'd13535 : data_rom <= {16'd31553, 16'd8839};
                15'd13536 : data_rom <= {16'd31554, 16'd8836};
                15'd13537 : data_rom <= {16'd31554, 16'd8833};
                15'd13538 : data_rom <= {16'd31555, 16'd8830};
                15'd13539 : data_rom <= {16'd31556, 16'd8827};
                15'd13540 : data_rom <= {16'd31557, 16'd8824};
                15'd13541 : data_rom <= {16'd31558, 16'd8821};
                15'd13542 : data_rom <= {16'd31559, 16'd8818};
                15'd13543 : data_rom <= {16'd31559, 16'd8815};
                15'd13544 : data_rom <= {16'd31560, 16'd8812};
                15'd13545 : data_rom <= {16'd31561, 16'd8809};
                15'd13546 : data_rom <= {16'd31562, 16'd8806};
                15'd13547 : data_rom <= {16'd31563, 16'd8803};
                15'd13548 : data_rom <= {16'd31564, 16'd8800};
                15'd13549 : data_rom <= {16'd31565, 16'd8797};
                15'd13550 : data_rom <= {16'd31565, 16'd8794};
                15'd13551 : data_rom <= {16'd31566, 16'd8791};
                15'd13552 : data_rom <= {16'd31567, 16'd8788};
                15'd13553 : data_rom <= {16'd31568, 16'd8785};
                15'd13554 : data_rom <= {16'd31569, 16'd8782};
                15'd13555 : data_rom <= {16'd31570, 16'd8779};
                15'd13556 : data_rom <= {16'd31570, 16'd8776};
                15'd13557 : data_rom <= {16'd31571, 16'd8772};
                15'd13558 : data_rom <= {16'd31572, 16'd8769};
                15'd13559 : data_rom <= {16'd31573, 16'd8766};
                15'd13560 : data_rom <= {16'd31574, 16'd8763};
                15'd13561 : data_rom <= {16'd31575, 16'd8760};
                15'd13562 : data_rom <= {16'd31575, 16'd8757};
                15'd13563 : data_rom <= {16'd31576, 16'd8754};
                15'd13564 : data_rom <= {16'd31577, 16'd8751};
                15'd13565 : data_rom <= {16'd31578, 16'd8748};
                15'd13566 : data_rom <= {16'd31579, 16'd8745};
                15'd13567 : data_rom <= {16'd31580, 16'd8742};
                15'd13568 : data_rom <= {16'd31581, 16'd8739};
                15'd13569 : data_rom <= {16'd31581, 16'd8736};
                15'd13570 : data_rom <= {16'd31582, 16'd8733};
                15'd13571 : data_rom <= {16'd31583, 16'd8730};
                15'd13572 : data_rom <= {16'd31584, 16'd8727};
                15'd13573 : data_rom <= {16'd31585, 16'd8724};
                15'd13574 : data_rom <= {16'd31586, 16'd8721};
                15'd13575 : data_rom <= {16'd31586, 16'd8718};
                15'd13576 : data_rom <= {16'd31587, 16'd8715};
                15'd13577 : data_rom <= {16'd31588, 16'd8712};
                15'd13578 : data_rom <= {16'd31589, 16'd8709};
                15'd13579 : data_rom <= {16'd31590, 16'd8706};
                15'd13580 : data_rom <= {16'd31591, 16'd8703};
                15'd13581 : data_rom <= {16'd31591, 16'd8700};
                15'd13582 : data_rom <= {16'd31592, 16'd8697};
                15'd13583 : data_rom <= {16'd31593, 16'd8694};
                15'd13584 : data_rom <= {16'd31594, 16'd8691};
                15'd13585 : data_rom <= {16'd31595, 16'd8688};
                15'd13586 : data_rom <= {16'd31596, 16'd8685};
                15'd13587 : data_rom <= {16'd31596, 16'd8682};
                15'd13588 : data_rom <= {16'd31597, 16'd8679};
                15'd13589 : data_rom <= {16'd31598, 16'd8676};
                15'd13590 : data_rom <= {16'd31599, 16'd8673};
                15'd13591 : data_rom <= {16'd31600, 16'd8670};
                15'd13592 : data_rom <= {16'd31601, 16'd8666};
                15'd13593 : data_rom <= {16'd31601, 16'd8663};
                15'd13594 : data_rom <= {16'd31602, 16'd8660};
                15'd13595 : data_rom <= {16'd31603, 16'd8657};
                15'd13596 : data_rom <= {16'd31604, 16'd8654};
                15'd13597 : data_rom <= {16'd31605, 16'd8651};
                15'd13598 : data_rom <= {16'd31606, 16'd8648};
                15'd13599 : data_rom <= {16'd31606, 16'd8645};
                15'd13600 : data_rom <= {16'd31607, 16'd8642};
                15'd13601 : data_rom <= {16'd31608, 16'd8639};
                15'd13602 : data_rom <= {16'd31609, 16'd8636};
                15'd13603 : data_rom <= {16'd31610, 16'd8633};
                15'd13604 : data_rom <= {16'd31610, 16'd8630};
                15'd13605 : data_rom <= {16'd31611, 16'd8627};
                15'd13606 : data_rom <= {16'd31612, 16'd8624};
                15'd13607 : data_rom <= {16'd31613, 16'd8621};
                15'd13608 : data_rom <= {16'd31614, 16'd8618};
                15'd13609 : data_rom <= {16'd31615, 16'd8615};
                15'd13610 : data_rom <= {16'd31615, 16'd8612};
                15'd13611 : data_rom <= {16'd31616, 16'd8609};
                15'd13612 : data_rom <= {16'd31617, 16'd8606};
                15'd13613 : data_rom <= {16'd31618, 16'd8603};
                15'd13614 : data_rom <= {16'd31619, 16'd8600};
                15'd13615 : data_rom <= {16'd31620, 16'd8597};
                15'd13616 : data_rom <= {16'd31620, 16'd8594};
                15'd13617 : data_rom <= {16'd31621, 16'd8591};
                15'd13618 : data_rom <= {16'd31622, 16'd8588};
                15'd13619 : data_rom <= {16'd31623, 16'd8585};
                15'd13620 : data_rom <= {16'd31624, 16'd8582};
                15'd13621 : data_rom <= {16'd31625, 16'd8579};
                15'd13622 : data_rom <= {16'd31625, 16'd8576};
                15'd13623 : data_rom <= {16'd31626, 16'd8573};
                15'd13624 : data_rom <= {16'd31627, 16'd8570};
                15'd13625 : data_rom <= {16'd31628, 16'd8566};
                15'd13626 : data_rom <= {16'd31629, 16'd8563};
                15'd13627 : data_rom <= {16'd31629, 16'd8560};
                15'd13628 : data_rom <= {16'd31630, 16'd8557};
                15'd13629 : data_rom <= {16'd31631, 16'd8554};
                15'd13630 : data_rom <= {16'd31632, 16'd8551};
                15'd13631 : data_rom <= {16'd31633, 16'd8548};
                15'd13632 : data_rom <= {16'd31634, 16'd8545};
                15'd13633 : data_rom <= {16'd31634, 16'd8542};
                15'd13634 : data_rom <= {16'd31635, 16'd8539};
                15'd13635 : data_rom <= {16'd31636, 16'd8536};
                15'd13636 : data_rom <= {16'd31637, 16'd8533};
                15'd13637 : data_rom <= {16'd31638, 16'd8530};
                15'd13638 : data_rom <= {16'd31638, 16'd8527};
                15'd13639 : data_rom <= {16'd31639, 16'd8524};
                15'd13640 : data_rom <= {16'd31640, 16'd8521};
                15'd13641 : data_rom <= {16'd31641, 16'd8518};
                15'd13642 : data_rom <= {16'd31642, 16'd8515};
                15'd13643 : data_rom <= {16'd31643, 16'd8512};
                15'd13644 : data_rom <= {16'd31643, 16'd8509};
                15'd13645 : data_rom <= {16'd31644, 16'd8506};
                15'd13646 : data_rom <= {16'd31645, 16'd8503};
                15'd13647 : data_rom <= {16'd31646, 16'd8500};
                15'd13648 : data_rom <= {16'd31647, 16'd8497};
                15'd13649 : data_rom <= {16'd31647, 16'd8494};
                15'd13650 : data_rom <= {16'd31648, 16'd8491};
                15'd13651 : data_rom <= {16'd31649, 16'd8488};
                15'd13652 : data_rom <= {16'd31650, 16'd8485};
                15'd13653 : data_rom <= {16'd31651, 16'd8482};
                15'd13654 : data_rom <= {16'd31651, 16'd8478};
                15'd13655 : data_rom <= {16'd31652, 16'd8475};
                15'd13656 : data_rom <= {16'd31653, 16'd8472};
                15'd13657 : data_rom <= {16'd31654, 16'd8469};
                15'd13658 : data_rom <= {16'd31655, 16'd8466};
                15'd13659 : data_rom <= {16'd31656, 16'd8463};
                15'd13660 : data_rom <= {16'd31656, 16'd8460};
                15'd13661 : data_rom <= {16'd31657, 16'd8457};
                15'd13662 : data_rom <= {16'd31658, 16'd8454};
                15'd13663 : data_rom <= {16'd31659, 16'd8451};
                15'd13664 : data_rom <= {16'd31660, 16'd8448};
                15'd13665 : data_rom <= {16'd31660, 16'd8445};
                15'd13666 : data_rom <= {16'd31661, 16'd8442};
                15'd13667 : data_rom <= {16'd31662, 16'd8439};
                15'd13668 : data_rom <= {16'd31663, 16'd8436};
                15'd13669 : data_rom <= {16'd31664, 16'd8433};
                15'd13670 : data_rom <= {16'd31664, 16'd8430};
                15'd13671 : data_rom <= {16'd31665, 16'd8427};
                15'd13672 : data_rom <= {16'd31666, 16'd8424};
                15'd13673 : data_rom <= {16'd31667, 16'd8421};
                15'd13674 : data_rom <= {16'd31668, 16'd8418};
                15'd13675 : data_rom <= {16'd31668, 16'd8415};
                15'd13676 : data_rom <= {16'd31669, 16'd8412};
                15'd13677 : data_rom <= {16'd31670, 16'd8409};
                15'd13678 : data_rom <= {16'd31671, 16'd8406};
                15'd13679 : data_rom <= {16'd31672, 16'd8403};
                15'd13680 : data_rom <= {16'd31673, 16'd8400};
                15'd13681 : data_rom <= {16'd31673, 16'd8397};
                15'd13682 : data_rom <= {16'd31674, 16'd8393};
                15'd13683 : data_rom <= {16'd31675, 16'd8390};
                15'd13684 : data_rom <= {16'd31676, 16'd8387};
                15'd13685 : data_rom <= {16'd31677, 16'd8384};
                15'd13686 : data_rom <= {16'd31677, 16'd8381};
                15'd13687 : data_rom <= {16'd31678, 16'd8378};
                15'd13688 : data_rom <= {16'd31679, 16'd8375};
                15'd13689 : data_rom <= {16'd31680, 16'd8372};
                15'd13690 : data_rom <= {16'd31681, 16'd8369};
                15'd13691 : data_rom <= {16'd31681, 16'd8366};
                15'd13692 : data_rom <= {16'd31682, 16'd8363};
                15'd13693 : data_rom <= {16'd31683, 16'd8360};
                15'd13694 : data_rom <= {16'd31684, 16'd8357};
                15'd13695 : data_rom <= {16'd31685, 16'd8354};
                15'd13696 : data_rom <= {16'd31685, 16'd8351};
                15'd13697 : data_rom <= {16'd31686, 16'd8348};
                15'd13698 : data_rom <= {16'd31687, 16'd8345};
                15'd13699 : data_rom <= {16'd31688, 16'd8342};
                15'd13700 : data_rom <= {16'd31689, 16'd8339};
                15'd13701 : data_rom <= {16'd31689, 16'd8336};
                15'd13702 : data_rom <= {16'd31690, 16'd8333};
                15'd13703 : data_rom <= {16'd31691, 16'd8330};
                15'd13704 : data_rom <= {16'd31692, 16'd8327};
                15'd13705 : data_rom <= {16'd31693, 16'd8324};
                15'd13706 : data_rom <= {16'd31693, 16'd8321};
                15'd13707 : data_rom <= {16'd31694, 16'd8318};
                15'd13708 : data_rom <= {16'd31695, 16'd8315};
                15'd13709 : data_rom <= {16'd31696, 16'd8311};
                15'd13710 : data_rom <= {16'd31697, 16'd8308};
                15'd13711 : data_rom <= {16'd31697, 16'd8305};
                15'd13712 : data_rom <= {16'd31698, 16'd8302};
                15'd13713 : data_rom <= {16'd31699, 16'd8299};
                15'd13714 : data_rom <= {16'd31700, 16'd8296};
                15'd13715 : data_rom <= {16'd31701, 16'd8293};
                15'd13716 : data_rom <= {16'd31701, 16'd8290};
                15'd13717 : data_rom <= {16'd31702, 16'd8287};
                15'd13718 : data_rom <= {16'd31703, 16'd8284};
                15'd13719 : data_rom <= {16'd31704, 16'd8281};
                15'd13720 : data_rom <= {16'd31705, 16'd8278};
                15'd13721 : data_rom <= {16'd31705, 16'd8275};
                15'd13722 : data_rom <= {16'd31706, 16'd8272};
                15'd13723 : data_rom <= {16'd31707, 16'd8269};
                15'd13724 : data_rom <= {16'd31708, 16'd8266};
                15'd13725 : data_rom <= {16'd31708, 16'd8263};
                15'd13726 : data_rom <= {16'd31709, 16'd8260};
                15'd13727 : data_rom <= {16'd31710, 16'd8257};
                15'd13728 : data_rom <= {16'd31711, 16'd8254};
                15'd13729 : data_rom <= {16'd31712, 16'd8251};
                15'd13730 : data_rom <= {16'd31712, 16'd8248};
                15'd13731 : data_rom <= {16'd31713, 16'd8245};
                15'd13732 : data_rom <= {16'd31714, 16'd8242};
                15'd13733 : data_rom <= {16'd31715, 16'd8239};
                15'd13734 : data_rom <= {16'd31716, 16'd8235};
                15'd13735 : data_rom <= {16'd31716, 16'd8232};
                15'd13736 : data_rom <= {16'd31717, 16'd8229};
                15'd13737 : data_rom <= {16'd31718, 16'd8226};
                15'd13738 : data_rom <= {16'd31719, 16'd8223};
                15'd13739 : data_rom <= {16'd31720, 16'd8220};
                15'd13740 : data_rom <= {16'd31720, 16'd8217};
                15'd13741 : data_rom <= {16'd31721, 16'd8214};
                15'd13742 : data_rom <= {16'd31722, 16'd8211};
                15'd13743 : data_rom <= {16'd31723, 16'd8208};
                15'd13744 : data_rom <= {16'd31723, 16'd8205};
                15'd13745 : data_rom <= {16'd31724, 16'd8202};
                15'd13746 : data_rom <= {16'd31725, 16'd8199};
                15'd13747 : data_rom <= {16'd31726, 16'd8196};
                15'd13748 : data_rom <= {16'd31727, 16'd8193};
                15'd13749 : data_rom <= {16'd31727, 16'd8190};
                15'd13750 : data_rom <= {16'd31728, 16'd8187};
                15'd13751 : data_rom <= {16'd31729, 16'd8184};
                15'd13752 : data_rom <= {16'd31730, 16'd8181};
                15'd13753 : data_rom <= {16'd31731, 16'd8178};
                15'd13754 : data_rom <= {16'd31731, 16'd8175};
                15'd13755 : data_rom <= {16'd31732, 16'd8172};
                15'd13756 : data_rom <= {16'd31733, 16'd8169};
                15'd13757 : data_rom <= {16'd31734, 16'd8166};
                15'd13758 : data_rom <= {16'd31734, 16'd8162};
                15'd13759 : data_rom <= {16'd31735, 16'd8159};
                15'd13760 : data_rom <= {16'd31736, 16'd8156};
                15'd13761 : data_rom <= {16'd31737, 16'd8153};
                15'd13762 : data_rom <= {16'd31738, 16'd8150};
                15'd13763 : data_rom <= {16'd31738, 16'd8147};
                15'd13764 : data_rom <= {16'd31739, 16'd8144};
                15'd13765 : data_rom <= {16'd31740, 16'd8141};
                15'd13766 : data_rom <= {16'd31741, 16'd8138};
                15'd13767 : data_rom <= {16'd31741, 16'd8135};
                15'd13768 : data_rom <= {16'd31742, 16'd8132};
                15'd13769 : data_rom <= {16'd31743, 16'd8129};
                15'd13770 : data_rom <= {16'd31744, 16'd8126};
                15'd13771 : data_rom <= {16'd31745, 16'd8123};
                15'd13772 : data_rom <= {16'd31745, 16'd8120};
                15'd13773 : data_rom <= {16'd31746, 16'd8117};
                15'd13774 : data_rom <= {16'd31747, 16'd8114};
                15'd13775 : data_rom <= {16'd31748, 16'd8111};
                15'd13776 : data_rom <= {16'd31748, 16'd8108};
                15'd13777 : data_rom <= {16'd31749, 16'd8105};
                15'd13778 : data_rom <= {16'd31750, 16'd8102};
                15'd13779 : data_rom <= {16'd31751, 16'd8099};
                15'd13780 : data_rom <= {16'd31752, 16'd8096};
                15'd13781 : data_rom <= {16'd31752, 16'd8092};
                15'd13782 : data_rom <= {16'd31753, 16'd8089};
                15'd13783 : data_rom <= {16'd31754, 16'd8086};
                15'd13784 : data_rom <= {16'd31755, 16'd8083};
                15'd13785 : data_rom <= {16'd31755, 16'd8080};
                15'd13786 : data_rom <= {16'd31756, 16'd8077};
                15'd13787 : data_rom <= {16'd31757, 16'd8074};
                15'd13788 : data_rom <= {16'd31758, 16'd8071};
                15'd13789 : data_rom <= {16'd31759, 16'd8068};
                15'd13790 : data_rom <= {16'd31759, 16'd8065};
                15'd13791 : data_rom <= {16'd31760, 16'd8062};
                15'd13792 : data_rom <= {16'd31761, 16'd8059};
                15'd13793 : data_rom <= {16'd31762, 16'd8056};
                15'd13794 : data_rom <= {16'd31762, 16'd8053};
                15'd13795 : data_rom <= {16'd31763, 16'd8050};
                15'd13796 : data_rom <= {16'd31764, 16'd8047};
                15'd13797 : data_rom <= {16'd31765, 16'd8044};
                15'd13798 : data_rom <= {16'd31766, 16'd8041};
                15'd13799 : data_rom <= {16'd31766, 16'd8038};
                15'd13800 : data_rom <= {16'd31767, 16'd8035};
                15'd13801 : data_rom <= {16'd31768, 16'd8032};
                15'd13802 : data_rom <= {16'd31769, 16'd8029};
                15'd13803 : data_rom <= {16'd31769, 16'd8025};
                15'd13804 : data_rom <= {16'd31770, 16'd8022};
                15'd13805 : data_rom <= {16'd31771, 16'd8019};
                15'd13806 : data_rom <= {16'd31772, 16'd8016};
                15'd13807 : data_rom <= {16'd31772, 16'd8013};
                15'd13808 : data_rom <= {16'd31773, 16'd8010};
                15'd13809 : data_rom <= {16'd31774, 16'd8007};
                15'd13810 : data_rom <= {16'd31775, 16'd8004};
                15'd13811 : data_rom <= {16'd31776, 16'd8001};
                15'd13812 : data_rom <= {16'd31776, 16'd7998};
                15'd13813 : data_rom <= {16'd31777, 16'd7995};
                15'd13814 : data_rom <= {16'd31778, 16'd7992};
                15'd13815 : data_rom <= {16'd31779, 16'd7989};
                15'd13816 : data_rom <= {16'd31779, 16'd7986};
                15'd13817 : data_rom <= {16'd31780, 16'd7983};
                15'd13818 : data_rom <= {16'd31781, 16'd7980};
                15'd13819 : data_rom <= {16'd31782, 16'd7977};
                15'd13820 : data_rom <= {16'd31782, 16'd7974};
                15'd13821 : data_rom <= {16'd31783, 16'd7971};
                15'd13822 : data_rom <= {16'd31784, 16'd7968};
                15'd13823 : data_rom <= {16'd31785, 16'd7965};
                15'd13824 : data_rom <= {16'd31785, 16'd7962};
                15'd13825 : data_rom <= {16'd31786, 16'd7958};
                15'd13826 : data_rom <= {16'd31787, 16'd7955};
                15'd13827 : data_rom <= {16'd31788, 16'd7952};
                15'd13828 : data_rom <= {16'd31789, 16'd7949};
                15'd13829 : data_rom <= {16'd31789, 16'd7946};
                15'd13830 : data_rom <= {16'd31790, 16'd7943};
                15'd13831 : data_rom <= {16'd31791, 16'd7940};
                15'd13832 : data_rom <= {16'd31792, 16'd7937};
                15'd13833 : data_rom <= {16'd31792, 16'd7934};
                15'd13834 : data_rom <= {16'd31793, 16'd7931};
                15'd13835 : data_rom <= {16'd31794, 16'd7928};
                15'd13836 : data_rom <= {16'd31795, 16'd7925};
                15'd13837 : data_rom <= {16'd31795, 16'd7922};
                15'd13838 : data_rom <= {16'd31796, 16'd7919};
                15'd13839 : data_rom <= {16'd31797, 16'd7916};
                15'd13840 : data_rom <= {16'd31798, 16'd7913};
                15'd13841 : data_rom <= {16'd31798, 16'd7910};
                15'd13842 : data_rom <= {16'd31799, 16'd7907};
                15'd13843 : data_rom <= {16'd31800, 16'd7904};
                15'd13844 : data_rom <= {16'd31801, 16'd7901};
                15'd13845 : data_rom <= {16'd31801, 16'd7898};
                15'd13846 : data_rom <= {16'd31802, 16'd7894};
                15'd13847 : data_rom <= {16'd31803, 16'd7891};
                15'd13848 : data_rom <= {16'd31804, 16'd7888};
                15'd13849 : data_rom <= {16'd31804, 16'd7885};
                15'd13850 : data_rom <= {16'd31805, 16'd7882};
                15'd13851 : data_rom <= {16'd31806, 16'd7879};
                15'd13852 : data_rom <= {16'd31807, 16'd7876};
                15'd13853 : data_rom <= {16'd31807, 16'd7873};
                15'd13854 : data_rom <= {16'd31808, 16'd7870};
                15'd13855 : data_rom <= {16'd31809, 16'd7867};
                15'd13856 : data_rom <= {16'd31810, 16'd7864};
                15'd13857 : data_rom <= {16'd31811, 16'd7861};
                15'd13858 : data_rom <= {16'd31811, 16'd7858};
                15'd13859 : data_rom <= {16'd31812, 16'd7855};
                15'd13860 : data_rom <= {16'd31813, 16'd7852};
                15'd13861 : data_rom <= {16'd31814, 16'd7849};
                15'd13862 : data_rom <= {16'd31814, 16'd7846};
                15'd13863 : data_rom <= {16'd31815, 16'd7843};
                15'd13864 : data_rom <= {16'd31816, 16'd7840};
                15'd13865 : data_rom <= {16'd31817, 16'd7837};
                15'd13866 : data_rom <= {16'd31817, 16'd7833};
                15'd13867 : data_rom <= {16'd31818, 16'd7830};
                15'd13868 : data_rom <= {16'd31819, 16'd7827};
                15'd13869 : data_rom <= {16'd31820, 16'd7824};
                15'd13870 : data_rom <= {16'd31820, 16'd7821};
                15'd13871 : data_rom <= {16'd31821, 16'd7818};
                15'd13872 : data_rom <= {16'd31822, 16'd7815};
                15'd13873 : data_rom <= {16'd31823, 16'd7812};
                15'd13874 : data_rom <= {16'd31823, 16'd7809};
                15'd13875 : data_rom <= {16'd31824, 16'd7806};
                15'd13876 : data_rom <= {16'd31825, 16'd7803};
                15'd13877 : data_rom <= {16'd31826, 16'd7800};
                15'd13878 : data_rom <= {16'd31826, 16'd7797};
                15'd13879 : data_rom <= {16'd31827, 16'd7794};
                15'd13880 : data_rom <= {16'd31828, 16'd7791};
                15'd13881 : data_rom <= {16'd31829, 16'd7788};
                15'd13882 : data_rom <= {16'd31829, 16'd7785};
                15'd13883 : data_rom <= {16'd31830, 16'd7782};
                15'd13884 : data_rom <= {16'd31831, 16'd7779};
                15'd13885 : data_rom <= {16'd31831, 16'd7775};
                15'd13886 : data_rom <= {16'd31832, 16'd7772};
                15'd13887 : data_rom <= {16'd31833, 16'd7769};
                15'd13888 : data_rom <= {16'd31834, 16'd7766};
                15'd13889 : data_rom <= {16'd31834, 16'd7763};
                15'd13890 : data_rom <= {16'd31835, 16'd7760};
                15'd13891 : data_rom <= {16'd31836, 16'd7757};
                15'd13892 : data_rom <= {16'd31837, 16'd7754};
                15'd13893 : data_rom <= {16'd31837, 16'd7751};
                15'd13894 : data_rom <= {16'd31838, 16'd7748};
                15'd13895 : data_rom <= {16'd31839, 16'd7745};
                15'd13896 : data_rom <= {16'd31840, 16'd7742};
                15'd13897 : data_rom <= {16'd31840, 16'd7739};
                15'd13898 : data_rom <= {16'd31841, 16'd7736};
                15'd13899 : data_rom <= {16'd31842, 16'd7733};
                15'd13900 : data_rom <= {16'd31843, 16'd7730};
                15'd13901 : data_rom <= {16'd31843, 16'd7727};
                15'd13902 : data_rom <= {16'd31844, 16'd7724};
                15'd13903 : data_rom <= {16'd31845, 16'd7721};
                15'd13904 : data_rom <= {16'd31846, 16'd7717};
                15'd13905 : data_rom <= {16'd31846, 16'd7714};
                15'd13906 : data_rom <= {16'd31847, 16'd7711};
                15'd13907 : data_rom <= {16'd31848, 16'd7708};
                15'd13908 : data_rom <= {16'd31849, 16'd7705};
                15'd13909 : data_rom <= {16'd31849, 16'd7702};
                15'd13910 : data_rom <= {16'd31850, 16'd7699};
                15'd13911 : data_rom <= {16'd31851, 16'd7696};
                15'd13912 : data_rom <= {16'd31852, 16'd7693};
                15'd13913 : data_rom <= {16'd31852, 16'd7690};
                15'd13914 : data_rom <= {16'd31853, 16'd7687};
                15'd13915 : data_rom <= {16'd31854, 16'd7684};
                15'd13916 : data_rom <= {16'd31854, 16'd7681};
                15'd13917 : data_rom <= {16'd31855, 16'd7678};
                15'd13918 : data_rom <= {16'd31856, 16'd7675};
                15'd13919 : data_rom <= {16'd31857, 16'd7672};
                15'd13920 : data_rom <= {16'd31857, 16'd7669};
                15'd13921 : data_rom <= {16'd31858, 16'd7666};
                15'd13922 : data_rom <= {16'd31859, 16'd7663};
                15'd13923 : data_rom <= {16'd31860, 16'd7659};
                15'd13924 : data_rom <= {16'd31860, 16'd7656};
                15'd13925 : data_rom <= {16'd31861, 16'd7653};
                15'd13926 : data_rom <= {16'd31862, 16'd7650};
                15'd13927 : data_rom <= {16'd31863, 16'd7647};
                15'd13928 : data_rom <= {16'd31863, 16'd7644};
                15'd13929 : data_rom <= {16'd31864, 16'd7641};
                15'd13930 : data_rom <= {16'd31865, 16'd7638};
                15'd13931 : data_rom <= {16'd31865, 16'd7635};
                15'd13932 : data_rom <= {16'd31866, 16'd7632};
                15'd13933 : data_rom <= {16'd31867, 16'd7629};
                15'd13934 : data_rom <= {16'd31868, 16'd7626};
                15'd13935 : data_rom <= {16'd31868, 16'd7623};
                15'd13936 : data_rom <= {16'd31869, 16'd7620};
                15'd13937 : data_rom <= {16'd31870, 16'd7617};
                15'd13938 : data_rom <= {16'd31871, 16'd7614};
                15'd13939 : data_rom <= {16'd31871, 16'd7611};
                15'd13940 : data_rom <= {16'd31872, 16'd7608};
                15'd13941 : data_rom <= {16'd31873, 16'd7604};
                15'd13942 : data_rom <= {16'd31874, 16'd7601};
                15'd13943 : data_rom <= {16'd31874, 16'd7598};
                15'd13944 : data_rom <= {16'd31875, 16'd7595};
                15'd13945 : data_rom <= {16'd31876, 16'd7592};
                15'd13946 : data_rom <= {16'd31876, 16'd7589};
                15'd13947 : data_rom <= {16'd31877, 16'd7586};
                15'd13948 : data_rom <= {16'd31878, 16'd7583};
                15'd13949 : data_rom <= {16'd31879, 16'd7580};
                15'd13950 : data_rom <= {16'd31879, 16'd7577};
                15'd13951 : data_rom <= {16'd31880, 16'd7574};
                15'd13952 : data_rom <= {16'd31881, 16'd7571};
                15'd13953 : data_rom <= {16'd31882, 16'd7568};
                15'd13954 : data_rom <= {16'd31882, 16'd7565};
                15'd13955 : data_rom <= {16'd31883, 16'd7562};
                15'd13956 : data_rom <= {16'd31884, 16'd7559};
                15'd13957 : data_rom <= {16'd31884, 16'd7556};
                15'd13958 : data_rom <= {16'd31885, 16'd7553};
                15'd13959 : data_rom <= {16'd31886, 16'd7549};
                15'd13960 : data_rom <= {16'd31887, 16'd7546};
                15'd13961 : data_rom <= {16'd31887, 16'd7543};
                15'd13962 : data_rom <= {16'd31888, 16'd7540};
                15'd13963 : data_rom <= {16'd31889, 16'd7537};
                15'd13964 : data_rom <= {16'd31889, 16'd7534};
                15'd13965 : data_rom <= {16'd31890, 16'd7531};
                15'd13966 : data_rom <= {16'd31891, 16'd7528};
                15'd13967 : data_rom <= {16'd31892, 16'd7525};
                15'd13968 : data_rom <= {16'd31892, 16'd7522};
                15'd13969 : data_rom <= {16'd31893, 16'd7519};
                15'd13970 : data_rom <= {16'd31894, 16'd7516};
                15'd13971 : data_rom <= {16'd31895, 16'd7513};
                15'd13972 : data_rom <= {16'd31895, 16'd7510};
                15'd13973 : data_rom <= {16'd31896, 16'd7507};
                15'd13974 : data_rom <= {16'd31897, 16'd7504};
                15'd13975 : data_rom <= {16'd31897, 16'd7501};
                15'd13976 : data_rom <= {16'd31898, 16'd7497};
                15'd13977 : data_rom <= {16'd31899, 16'd7494};
                15'd13978 : data_rom <= {16'd31900, 16'd7491};
                15'd13979 : data_rom <= {16'd31900, 16'd7488};
                15'd13980 : data_rom <= {16'd31901, 16'd7485};
                15'd13981 : data_rom <= {16'd31902, 16'd7482};
                15'd13982 : data_rom <= {16'd31902, 16'd7479};
                15'd13983 : data_rom <= {16'd31903, 16'd7476};
                15'd13984 : data_rom <= {16'd31904, 16'd7473};
                15'd13985 : data_rom <= {16'd31905, 16'd7470};
                15'd13986 : data_rom <= {16'd31905, 16'd7467};
                15'd13987 : data_rom <= {16'd31906, 16'd7464};
                15'd13988 : data_rom <= {16'd31907, 16'd7461};
                15'd13989 : data_rom <= {16'd31907, 16'd7458};
                15'd13990 : data_rom <= {16'd31908, 16'd7455};
                15'd13991 : data_rom <= {16'd31909, 16'd7452};
                15'd13992 : data_rom <= {16'd31910, 16'd7449};
                15'd13993 : data_rom <= {16'd31910, 16'd7445};
                15'd13994 : data_rom <= {16'd31911, 16'd7442};
                15'd13995 : data_rom <= {16'd31912, 16'd7439};
                15'd13996 : data_rom <= {16'd31912, 16'd7436};
                15'd13997 : data_rom <= {16'd31913, 16'd7433};
                15'd13998 : data_rom <= {16'd31914, 16'd7430};
                15'd13999 : data_rom <= {16'd31915, 16'd7427};
                15'd14000 : data_rom <= {16'd31915, 16'd7424};
                15'd14001 : data_rom <= {16'd31916, 16'd7421};
                15'd14002 : data_rom <= {16'd31917, 16'd7418};
                15'd14003 : data_rom <= {16'd31917, 16'd7415};
                15'd14004 : data_rom <= {16'd31918, 16'd7412};
                15'd14005 : data_rom <= {16'd31919, 16'd7409};
                15'd14006 : data_rom <= {16'd31920, 16'd7406};
                15'd14007 : data_rom <= {16'd31920, 16'd7403};
                15'd14008 : data_rom <= {16'd31921, 16'd7400};
                15'd14009 : data_rom <= {16'd31922, 16'd7397};
                15'd14010 : data_rom <= {16'd31922, 16'd7393};
                15'd14011 : data_rom <= {16'd31923, 16'd7390};
                15'd14012 : data_rom <= {16'd31924, 16'd7387};
                15'd14013 : data_rom <= {16'd31925, 16'd7384};
                15'd14014 : data_rom <= {16'd31925, 16'd7381};
                15'd14015 : data_rom <= {16'd31926, 16'd7378};
                15'd14016 : data_rom <= {16'd31927, 16'd7375};
                15'd14017 : data_rom <= {16'd31927, 16'd7372};
                15'd14018 : data_rom <= {16'd31928, 16'd7369};
                15'd14019 : data_rom <= {16'd31929, 16'd7366};
                15'd14020 : data_rom <= {16'd31929, 16'd7363};
                15'd14021 : data_rom <= {16'd31930, 16'd7360};
                15'd14022 : data_rom <= {16'd31931, 16'd7357};
                15'd14023 : data_rom <= {16'd31932, 16'd7354};
                15'd14024 : data_rom <= {16'd31932, 16'd7351};
                15'd14025 : data_rom <= {16'd31933, 16'd7348};
                15'd14026 : data_rom <= {16'd31934, 16'd7344};
                15'd14027 : data_rom <= {16'd31934, 16'd7341};
                15'd14028 : data_rom <= {16'd31935, 16'd7338};
                15'd14029 : data_rom <= {16'd31936, 16'd7335};
                15'd14030 : data_rom <= {16'd31937, 16'd7332};
                15'd14031 : data_rom <= {16'd31937, 16'd7329};
                15'd14032 : data_rom <= {16'd31938, 16'd7326};
                15'd14033 : data_rom <= {16'd31939, 16'd7323};
                15'd14034 : data_rom <= {16'd31939, 16'd7320};
                15'd14035 : data_rom <= {16'd31940, 16'd7317};
                15'd14036 : data_rom <= {16'd31941, 16'd7314};
                15'd14037 : data_rom <= {16'd31941, 16'd7311};
                15'd14038 : data_rom <= {16'd31942, 16'd7308};
                15'd14039 : data_rom <= {16'd31943, 16'd7305};
                15'd14040 : data_rom <= {16'd31944, 16'd7302};
                15'd14041 : data_rom <= {16'd31944, 16'd7299};
                15'd14042 : data_rom <= {16'd31945, 16'd7295};
                15'd14043 : data_rom <= {16'd31946, 16'd7292};
                15'd14044 : data_rom <= {16'd31946, 16'd7289};
                15'd14045 : data_rom <= {16'd31947, 16'd7286};
                15'd14046 : data_rom <= {16'd31948, 16'd7283};
                15'd14047 : data_rom <= {16'd31948, 16'd7280};
                15'd14048 : data_rom <= {16'd31949, 16'd7277};
                15'd14049 : data_rom <= {16'd31950, 16'd7274};
                15'd14050 : data_rom <= {16'd31951, 16'd7271};
                15'd14051 : data_rom <= {16'd31951, 16'd7268};
                15'd14052 : data_rom <= {16'd31952, 16'd7265};
                15'd14053 : data_rom <= {16'd31953, 16'd7262};
                15'd14054 : data_rom <= {16'd31953, 16'd7259};
                15'd14055 : data_rom <= {16'd31954, 16'd7256};
                15'd14056 : data_rom <= {16'd31955, 16'd7253};
                15'd14057 : data_rom <= {16'd31955, 16'd7250};
                15'd14058 : data_rom <= {16'd31956, 16'd7246};
                15'd14059 : data_rom <= {16'd31957, 16'd7243};
                15'd14060 : data_rom <= {16'd31957, 16'd7240};
                15'd14061 : data_rom <= {16'd31958, 16'd7237};
                15'd14062 : data_rom <= {16'd31959, 16'd7234};
                15'd14063 : data_rom <= {16'd31960, 16'd7231};
                15'd14064 : data_rom <= {16'd31960, 16'd7228};
                15'd14065 : data_rom <= {16'd31961, 16'd7225};
                15'd14066 : data_rom <= {16'd31962, 16'd7222};
                15'd14067 : data_rom <= {16'd31962, 16'd7219};
                15'd14068 : data_rom <= {16'd31963, 16'd7216};
                15'd14069 : data_rom <= {16'd31964, 16'd7213};
                15'd14070 : data_rom <= {16'd31964, 16'd7210};
                15'd14071 : data_rom <= {16'd31965, 16'd7207};
                15'd14072 : data_rom <= {16'd31966, 16'd7204};
                15'd14073 : data_rom <= {16'd31966, 16'd7201};
                15'd14074 : data_rom <= {16'd31967, 16'd7197};
                15'd14075 : data_rom <= {16'd31968, 16'd7194};
                15'd14076 : data_rom <= {16'd31969, 16'd7191};
                15'd14077 : data_rom <= {16'd31969, 16'd7188};
                15'd14078 : data_rom <= {16'd31970, 16'd7185};
                15'd14079 : data_rom <= {16'd31971, 16'd7182};
                15'd14080 : data_rom <= {16'd31971, 16'd7179};
                15'd14081 : data_rom <= {16'd31972, 16'd7176};
                15'd14082 : data_rom <= {16'd31973, 16'd7173};
                15'd14083 : data_rom <= {16'd31973, 16'd7170};
                15'd14084 : data_rom <= {16'd31974, 16'd7167};
                15'd14085 : data_rom <= {16'd31975, 16'd7164};
                15'd14086 : data_rom <= {16'd31975, 16'd7161};
                15'd14087 : data_rom <= {16'd31976, 16'd7158};
                15'd14088 : data_rom <= {16'd31977, 16'd7155};
                15'd14089 : data_rom <= {16'd31977, 16'd7151};
                15'd14090 : data_rom <= {16'd31978, 16'd7148};
                15'd14091 : data_rom <= {16'd31979, 16'd7145};
                15'd14092 : data_rom <= {16'd31980, 16'd7142};
                15'd14093 : data_rom <= {16'd31980, 16'd7139};
                15'd14094 : data_rom <= {16'd31981, 16'd7136};
                15'd14095 : data_rom <= {16'd31982, 16'd7133};
                15'd14096 : data_rom <= {16'd31982, 16'd7130};
                15'd14097 : data_rom <= {16'd31983, 16'd7127};
                15'd14098 : data_rom <= {16'd31984, 16'd7124};
                15'd14099 : data_rom <= {16'd31984, 16'd7121};
                15'd14100 : data_rom <= {16'd31985, 16'd7118};
                15'd14101 : data_rom <= {16'd31986, 16'd7115};
                15'd14102 : data_rom <= {16'd31986, 16'd7112};
                15'd14103 : data_rom <= {16'd31987, 16'd7109};
                15'd14104 : data_rom <= {16'd31988, 16'd7105};
                15'd14105 : data_rom <= {16'd31988, 16'd7102};
                15'd14106 : data_rom <= {16'd31989, 16'd7099};
                15'd14107 : data_rom <= {16'd31990, 16'd7096};
                15'd14108 : data_rom <= {16'd31990, 16'd7093};
                15'd14109 : data_rom <= {16'd31991, 16'd7090};
                15'd14110 : data_rom <= {16'd31992, 16'd7087};
                15'd14111 : data_rom <= {16'd31992, 16'd7084};
                15'd14112 : data_rom <= {16'd31993, 16'd7081};
                15'd14113 : data_rom <= {16'd31994, 16'd7078};
                15'd14114 : data_rom <= {16'd31995, 16'd7075};
                15'd14115 : data_rom <= {16'd31995, 16'd7072};
                15'd14116 : data_rom <= {16'd31996, 16'd7069};
                15'd14117 : data_rom <= {16'd31997, 16'd7066};
                15'd14118 : data_rom <= {16'd31997, 16'd7063};
                15'd14119 : data_rom <= {16'd31998, 16'd7059};
                15'd14120 : data_rom <= {16'd31999, 16'd7056};
                15'd14121 : data_rom <= {16'd31999, 16'd7053};
                15'd14122 : data_rom <= {16'd32000, 16'd7050};
                15'd14123 : data_rom <= {16'd32001, 16'd7047};
                15'd14124 : data_rom <= {16'd32001, 16'd7044};
                15'd14125 : data_rom <= {16'd32002, 16'd7041};
                15'd14126 : data_rom <= {16'd32003, 16'd7038};
                15'd14127 : data_rom <= {16'd32003, 16'd7035};
                15'd14128 : data_rom <= {16'd32004, 16'd7032};
                15'd14129 : data_rom <= {16'd32005, 16'd7029};
                15'd14130 : data_rom <= {16'd32005, 16'd7026};
                15'd14131 : data_rom <= {16'd32006, 16'd7023};
                15'd14132 : data_rom <= {16'd32007, 16'd7020};
                15'd14133 : data_rom <= {16'd32007, 16'd7016};
                15'd14134 : data_rom <= {16'd32008, 16'd7013};
                15'd14135 : data_rom <= {16'd32009, 16'd7010};
                15'd14136 : data_rom <= {16'd32009, 16'd7007};
                15'd14137 : data_rom <= {16'd32010, 16'd7004};
                15'd14138 : data_rom <= {16'd32011, 16'd7001};
                15'd14139 : data_rom <= {16'd32011, 16'd6998};
                15'd14140 : data_rom <= {16'd32012, 16'd6995};
                15'd14141 : data_rom <= {16'd32013, 16'd6992};
                15'd14142 : data_rom <= {16'd32013, 16'd6989};
                15'd14143 : data_rom <= {16'd32014, 16'd6986};
                15'd14144 : data_rom <= {16'd32015, 16'd6983};
                15'd14145 : data_rom <= {16'd32015, 16'd6980};
                15'd14146 : data_rom <= {16'd32016, 16'd6977};
                15'd14147 : data_rom <= {16'd32017, 16'd6974};
                15'd14148 : data_rom <= {16'd32017, 16'd6970};
                15'd14149 : data_rom <= {16'd32018, 16'd6967};
                15'd14150 : data_rom <= {16'd32019, 16'd6964};
                15'd14151 : data_rom <= {16'd32019, 16'd6961};
                15'd14152 : data_rom <= {16'd32020, 16'd6958};
                15'd14153 : data_rom <= {16'd32021, 16'd6955};
                15'd14154 : data_rom <= {16'd32021, 16'd6952};
                15'd14155 : data_rom <= {16'd32022, 16'd6949};
                15'd14156 : data_rom <= {16'd32023, 16'd6946};
                15'd14157 : data_rom <= {16'd32023, 16'd6943};
                15'd14158 : data_rom <= {16'd32024, 16'd6940};
                15'd14159 : data_rom <= {16'd32025, 16'd6937};
                15'd14160 : data_rom <= {16'd32025, 16'd6934};
                15'd14161 : data_rom <= {16'd32026, 16'd6931};
                15'd14162 : data_rom <= {16'd32027, 16'd6927};
                15'd14163 : data_rom <= {16'd32027, 16'd6924};
                15'd14164 : data_rom <= {16'd32028, 16'd6921};
                15'd14165 : data_rom <= {16'd32029, 16'd6918};
                15'd14166 : data_rom <= {16'd32029, 16'd6915};
                15'd14167 : data_rom <= {16'd32030, 16'd6912};
                15'd14168 : data_rom <= {16'd32031, 16'd6909};
                15'd14169 : data_rom <= {16'd32031, 16'd6906};
                15'd14170 : data_rom <= {16'd32032, 16'd6903};
                15'd14171 : data_rom <= {16'd32033, 16'd6900};
                15'd14172 : data_rom <= {16'd32033, 16'd6897};
                15'd14173 : data_rom <= {16'd32034, 16'd6894};
                15'd14174 : data_rom <= {16'd32035, 16'd6891};
                15'd14175 : data_rom <= {16'd32035, 16'd6888};
                15'd14176 : data_rom <= {16'd32036, 16'd6884};
                15'd14177 : data_rom <= {16'd32037, 16'd6881};
                15'd14178 : data_rom <= {16'd32037, 16'd6878};
                15'd14179 : data_rom <= {16'd32038, 16'd6875};
                15'd14180 : data_rom <= {16'd32039, 16'd6872};
                15'd14181 : data_rom <= {16'd32039, 16'd6869};
                15'd14182 : data_rom <= {16'd32040, 16'd6866};
                15'd14183 : data_rom <= {16'd32041, 16'd6863};
                15'd14184 : data_rom <= {16'd32041, 16'd6860};
                15'd14185 : data_rom <= {16'd32042, 16'd6857};
                15'd14186 : data_rom <= {16'd32043, 16'd6854};
                15'd14187 : data_rom <= {16'd32043, 16'd6851};
                15'd14188 : data_rom <= {16'd32044, 16'd6848};
                15'd14189 : data_rom <= {16'd32045, 16'd6845};
                15'd14190 : data_rom <= {16'd32045, 16'd6841};
                15'd14191 : data_rom <= {16'd32046, 16'd6838};
                15'd14192 : data_rom <= {16'd32047, 16'd6835};
                15'd14193 : data_rom <= {16'd32047, 16'd6832};
                15'd14194 : data_rom <= {16'd32048, 16'd6829};
                15'd14195 : data_rom <= {16'd32049, 16'd6826};
                15'd14196 : data_rom <= {16'd32049, 16'd6823};
                15'd14197 : data_rom <= {16'd32050, 16'd6820};
                15'd14198 : data_rom <= {16'd32050, 16'd6817};
                15'd14199 : data_rom <= {16'd32051, 16'd6814};
                15'd14200 : data_rom <= {16'd32052, 16'd6811};
                15'd14201 : data_rom <= {16'd32052, 16'd6808};
                15'd14202 : data_rom <= {16'd32053, 16'd6805};
                15'd14203 : data_rom <= {16'd32054, 16'd6802};
                15'd14204 : data_rom <= {16'd32054, 16'd6798};
                15'd14205 : data_rom <= {16'd32055, 16'd6795};
                15'd14206 : data_rom <= {16'd32056, 16'd6792};
                15'd14207 : data_rom <= {16'd32056, 16'd6789};
                15'd14208 : data_rom <= {16'd32057, 16'd6786};
                15'd14209 : data_rom <= {16'd32058, 16'd6783};
                15'd14210 : data_rom <= {16'd32058, 16'd6780};
                15'd14211 : data_rom <= {16'd32059, 16'd6777};
                15'd14212 : data_rom <= {16'd32060, 16'd6774};
                15'd14213 : data_rom <= {16'd32060, 16'd6771};
                15'd14214 : data_rom <= {16'd32061, 16'd6768};
                15'd14215 : data_rom <= {16'd32062, 16'd6765};
                15'd14216 : data_rom <= {16'd32062, 16'd6762};
                15'd14217 : data_rom <= {16'd32063, 16'd6759};
                15'd14218 : data_rom <= {16'd32063, 16'd6755};
                15'd14219 : data_rom <= {16'd32064, 16'd6752};
                15'd14220 : data_rom <= {16'd32065, 16'd6749};
                15'd14221 : data_rom <= {16'd32065, 16'd6746};
                15'd14222 : data_rom <= {16'd32066, 16'd6743};
                15'd14223 : data_rom <= {16'd32067, 16'd6740};
                15'd14224 : data_rom <= {16'd32067, 16'd6737};
                15'd14225 : data_rom <= {16'd32068, 16'd6734};
                15'd14226 : data_rom <= {16'd32069, 16'd6731};
                15'd14227 : data_rom <= {16'd32069, 16'd6728};
                15'd14228 : data_rom <= {16'd32070, 16'd6725};
                15'd14229 : data_rom <= {16'd32071, 16'd6722};
                15'd14230 : data_rom <= {16'd32071, 16'd6719};
                15'd14231 : data_rom <= {16'd32072, 16'd6715};
                15'd14232 : data_rom <= {16'd32073, 16'd6712};
                15'd14233 : data_rom <= {16'd32073, 16'd6709};
                15'd14234 : data_rom <= {16'd32074, 16'd6706};
                15'd14235 : data_rom <= {16'd32074, 16'd6703};
                15'd14236 : data_rom <= {16'd32075, 16'd6700};
                15'd14237 : data_rom <= {16'd32076, 16'd6697};
                15'd14238 : data_rom <= {16'd32076, 16'd6694};
                15'd14239 : data_rom <= {16'd32077, 16'd6691};
                15'd14240 : data_rom <= {16'd32078, 16'd6688};
                15'd14241 : data_rom <= {16'd32078, 16'd6685};
                15'd14242 : data_rom <= {16'd32079, 16'd6682};
                15'd14243 : data_rom <= {16'd32080, 16'd6679};
                15'd14244 : data_rom <= {16'd32080, 16'd6675};
                15'd14245 : data_rom <= {16'd32081, 16'd6672};
                15'd14246 : data_rom <= {16'd32082, 16'd6669};
                15'd14247 : data_rom <= {16'd32082, 16'd6666};
                15'd14248 : data_rom <= {16'd32083, 16'd6663};
                15'd14249 : data_rom <= {16'd32083, 16'd6660};
                15'd14250 : data_rom <= {16'd32084, 16'd6657};
                15'd14251 : data_rom <= {16'd32085, 16'd6654};
                15'd14252 : data_rom <= {16'd32085, 16'd6651};
                15'd14253 : data_rom <= {16'd32086, 16'd6648};
                15'd14254 : data_rom <= {16'd32087, 16'd6645};
                15'd14255 : data_rom <= {16'd32087, 16'd6642};
                15'd14256 : data_rom <= {16'd32088, 16'd6639};
                15'd14257 : data_rom <= {16'd32089, 16'd6635};
                15'd14258 : data_rom <= {16'd32089, 16'd6632};
                15'd14259 : data_rom <= {16'd32090, 16'd6629};
                15'd14260 : data_rom <= {16'd32090, 16'd6626};
                15'd14261 : data_rom <= {16'd32091, 16'd6623};
                15'd14262 : data_rom <= {16'd32092, 16'd6620};
                15'd14263 : data_rom <= {16'd32092, 16'd6617};
                15'd14264 : data_rom <= {16'd32093, 16'd6614};
                15'd14265 : data_rom <= {16'd32094, 16'd6611};
                15'd14266 : data_rom <= {16'd32094, 16'd6608};
                15'd14267 : data_rom <= {16'd32095, 16'd6605};
                15'd14268 : data_rom <= {16'd32096, 16'd6602};
                15'd14269 : data_rom <= {16'd32096, 16'd6599};
                15'd14270 : data_rom <= {16'd32097, 16'd6595};
                15'd14271 : data_rom <= {16'd32097, 16'd6592};
                15'd14272 : data_rom <= {16'd32098, 16'd6589};
                15'd14273 : data_rom <= {16'd32099, 16'd6586};
                15'd14274 : data_rom <= {16'd32099, 16'd6583};
                15'd14275 : data_rom <= {16'd32100, 16'd6580};
                15'd14276 : data_rom <= {16'd32101, 16'd6577};
                15'd14277 : data_rom <= {16'd32101, 16'd6574};
                15'd14278 : data_rom <= {16'd32102, 16'd6571};
                15'd14279 : data_rom <= {16'd32102, 16'd6568};
                15'd14280 : data_rom <= {16'd32103, 16'd6565};
                15'd14281 : data_rom <= {16'd32104, 16'd6562};
                15'd14282 : data_rom <= {16'd32104, 16'd6559};
                15'd14283 : data_rom <= {16'd32105, 16'd6555};
                15'd14284 : data_rom <= {16'd32106, 16'd6552};
                15'd14285 : data_rom <= {16'd32106, 16'd6549};
                15'd14286 : data_rom <= {16'd32107, 16'd6546};
                15'd14287 : data_rom <= {16'd32107, 16'd6543};
                15'd14288 : data_rom <= {16'd32108, 16'd6540};
                15'd14289 : data_rom <= {16'd32109, 16'd6537};
                15'd14290 : data_rom <= {16'd32109, 16'd6534};
                15'd14291 : data_rom <= {16'd32110, 16'd6531};
                15'd14292 : data_rom <= {16'd32111, 16'd6528};
                15'd14293 : data_rom <= {16'd32111, 16'd6525};
                15'd14294 : data_rom <= {16'd32112, 16'd6522};
                15'd14295 : data_rom <= {16'd32112, 16'd6519};
                15'd14296 : data_rom <= {16'd32113, 16'd6515};
                15'd14297 : data_rom <= {16'd32114, 16'd6512};
                15'd14298 : data_rom <= {16'd32114, 16'd6509};
                15'd14299 : data_rom <= {16'd32115, 16'd6506};
                15'd14300 : data_rom <= {16'd32116, 16'd6503};
                15'd14301 : data_rom <= {16'd32116, 16'd6500};
                15'd14302 : data_rom <= {16'd32117, 16'd6497};
                15'd14303 : data_rom <= {16'd32117, 16'd6494};
                15'd14304 : data_rom <= {16'd32118, 16'd6491};
                15'd14305 : data_rom <= {16'd32119, 16'd6488};
                15'd14306 : data_rom <= {16'd32119, 16'd6485};
                15'd14307 : data_rom <= {16'd32120, 16'd6482};
                15'd14308 : data_rom <= {16'd32121, 16'd6479};
                15'd14309 : data_rom <= {16'd32121, 16'd6475};
                15'd14310 : data_rom <= {16'd32122, 16'd6472};
                15'd14311 : data_rom <= {16'd32122, 16'd6469};
                15'd14312 : data_rom <= {16'd32123, 16'd6466};
                15'd14313 : data_rom <= {16'd32124, 16'd6463};
                15'd14314 : data_rom <= {16'd32124, 16'd6460};
                15'd14315 : data_rom <= {16'd32125, 16'd6457};
                15'd14316 : data_rom <= {16'd32126, 16'd6454};
                15'd14317 : data_rom <= {16'd32126, 16'd6451};
                15'd14318 : data_rom <= {16'd32127, 16'd6448};
                15'd14319 : data_rom <= {16'd32127, 16'd6445};
                15'd14320 : data_rom <= {16'd32128, 16'd6442};
                15'd14321 : data_rom <= {16'd32129, 16'd6438};
                15'd14322 : data_rom <= {16'd32129, 16'd6435};
                15'd14323 : data_rom <= {16'd32130, 16'd6432};
                15'd14324 : data_rom <= {16'd32130, 16'd6429};
                15'd14325 : data_rom <= {16'd32131, 16'd6426};
                15'd14326 : data_rom <= {16'd32132, 16'd6423};
                15'd14327 : data_rom <= {16'd32132, 16'd6420};
                15'd14328 : data_rom <= {16'd32133, 16'd6417};
                15'd14329 : data_rom <= {16'd32134, 16'd6414};
                15'd14330 : data_rom <= {16'd32134, 16'd6411};
                15'd14331 : data_rom <= {16'd32135, 16'd6408};
                15'd14332 : data_rom <= {16'd32135, 16'd6405};
                15'd14333 : data_rom <= {16'd32136, 16'd6402};
                15'd14334 : data_rom <= {16'd32137, 16'd6398};
                15'd14335 : data_rom <= {16'd32137, 16'd6395};
                15'd14336 : data_rom <= {16'd32138, 16'd6392};
                15'd14337 : data_rom <= {16'd32138, 16'd6389};
                15'd14338 : data_rom <= {16'd32139, 16'd6386};
                15'd14339 : data_rom <= {16'd32140, 16'd6383};
                15'd14340 : data_rom <= {16'd32140, 16'd6380};
                15'd14341 : data_rom <= {16'd32141, 16'd6377};
                15'd14342 : data_rom <= {16'd32142, 16'd6374};
                15'd14343 : data_rom <= {16'd32142, 16'd6371};
                15'd14344 : data_rom <= {16'd32143, 16'd6368};
                15'd14345 : data_rom <= {16'd32143, 16'd6365};
                15'd14346 : data_rom <= {16'd32144, 16'd6361};
                15'd14347 : data_rom <= {16'd32145, 16'd6358};
                15'd14348 : data_rom <= {16'd32145, 16'd6355};
                15'd14349 : data_rom <= {16'd32146, 16'd6352};
                15'd14350 : data_rom <= {16'd32146, 16'd6349};
                15'd14351 : data_rom <= {16'd32147, 16'd6346};
                15'd14352 : data_rom <= {16'd32148, 16'd6343};
                15'd14353 : data_rom <= {16'd32148, 16'd6340};
                15'd14354 : data_rom <= {16'd32149, 16'd6337};
                15'd14355 : data_rom <= {16'd32149, 16'd6334};
                15'd14356 : data_rom <= {16'd32150, 16'd6331};
                15'd14357 : data_rom <= {16'd32151, 16'd6328};
                15'd14358 : data_rom <= {16'd32151, 16'd6324};
                15'd14359 : data_rom <= {16'd32152, 16'd6321};
                15'd14360 : data_rom <= {16'd32152, 16'd6318};
                15'd14361 : data_rom <= {16'd32153, 16'd6315};
                15'd14362 : data_rom <= {16'd32154, 16'd6312};
                15'd14363 : data_rom <= {16'd32154, 16'd6309};
                15'd14364 : data_rom <= {16'd32155, 16'd6306};
                15'd14365 : data_rom <= {16'd32156, 16'd6303};
                15'd14366 : data_rom <= {16'd32156, 16'd6300};
                15'd14367 : data_rom <= {16'd32157, 16'd6297};
                15'd14368 : data_rom <= {16'd32157, 16'd6294};
                15'd14369 : data_rom <= {16'd32158, 16'd6291};
                15'd14370 : data_rom <= {16'd32159, 16'd6287};
                15'd14371 : data_rom <= {16'd32159, 16'd6284};
                15'd14372 : data_rom <= {16'd32160, 16'd6281};
                15'd14373 : data_rom <= {16'd32160, 16'd6278};
                15'd14374 : data_rom <= {16'd32161, 16'd6275};
                15'd14375 : data_rom <= {16'd32162, 16'd6272};
                15'd14376 : data_rom <= {16'd32162, 16'd6269};
                15'd14377 : data_rom <= {16'd32163, 16'd6266};
                15'd14378 : data_rom <= {16'd32163, 16'd6263};
                15'd14379 : data_rom <= {16'd32164, 16'd6260};
                15'd14380 : data_rom <= {16'd32165, 16'd6257};
                15'd14381 : data_rom <= {16'd32165, 16'd6254};
                15'd14382 : data_rom <= {16'd32166, 16'd6250};
                15'd14383 : data_rom <= {16'd32166, 16'd6247};
                15'd14384 : data_rom <= {16'd32167, 16'd6244};
                15'd14385 : data_rom <= {16'd32168, 16'd6241};
                15'd14386 : data_rom <= {16'd32168, 16'd6238};
                15'd14387 : data_rom <= {16'd32169, 16'd6235};
                15'd14388 : data_rom <= {16'd32169, 16'd6232};
                15'd14389 : data_rom <= {16'd32170, 16'd6229};
                15'd14390 : data_rom <= {16'd32171, 16'd6226};
                15'd14391 : data_rom <= {16'd32171, 16'd6223};
                15'd14392 : data_rom <= {16'd32172, 16'd6220};
                15'd14393 : data_rom <= {16'd32172, 16'd6217};
                15'd14394 : data_rom <= {16'd32173, 16'd6213};
                15'd14395 : data_rom <= {16'd32174, 16'd6210};
                15'd14396 : data_rom <= {16'd32174, 16'd6207};
                15'd14397 : data_rom <= {16'd32175, 16'd6204};
                15'd14398 : data_rom <= {16'd32175, 16'd6201};
                15'd14399 : data_rom <= {16'd32176, 16'd6198};
                15'd14400 : data_rom <= {16'd32176, 16'd6195};
                15'd14401 : data_rom <= {16'd32177, 16'd6192};
                15'd14402 : data_rom <= {16'd32178, 16'd6189};
                15'd14403 : data_rom <= {16'd32178, 16'd6186};
                15'd14404 : data_rom <= {16'd32179, 16'd6183};
                15'd14405 : data_rom <= {16'd32179, 16'd6180};
                15'd14406 : data_rom <= {16'd32180, 16'd6176};
                15'd14407 : data_rom <= {16'd32181, 16'd6173};
                15'd14408 : data_rom <= {16'd32181, 16'd6170};
                15'd14409 : data_rom <= {16'd32182, 16'd6167};
                15'd14410 : data_rom <= {16'd32182, 16'd6164};
                15'd14411 : data_rom <= {16'd32183, 16'd6161};
                15'd14412 : data_rom <= {16'd32184, 16'd6158};
                15'd14413 : data_rom <= {16'd32184, 16'd6155};
                15'd14414 : data_rom <= {16'd32185, 16'd6152};
                15'd14415 : data_rom <= {16'd32185, 16'd6149};
                15'd14416 : data_rom <= {16'd32186, 16'd6146};
                15'd14417 : data_rom <= {16'd32187, 16'd6142};
                15'd14418 : data_rom <= {16'd32187, 16'd6139};
                15'd14419 : data_rom <= {16'd32188, 16'd6136};
                15'd14420 : data_rom <= {16'd32188, 16'd6133};
                15'd14421 : data_rom <= {16'd32189, 16'd6130};
                15'd14422 : data_rom <= {16'd32189, 16'd6127};
                15'd14423 : data_rom <= {16'd32190, 16'd6124};
                15'd14424 : data_rom <= {16'd32191, 16'd6121};
                15'd14425 : data_rom <= {16'd32191, 16'd6118};
                15'd14426 : data_rom <= {16'd32192, 16'd6115};
                15'd14427 : data_rom <= {16'd32192, 16'd6112};
                15'd14428 : data_rom <= {16'd32193, 16'd6109};
                15'd14429 : data_rom <= {16'd32194, 16'd6105};
                15'd14430 : data_rom <= {16'd32194, 16'd6102};
                15'd14431 : data_rom <= {16'd32195, 16'd6099};
                15'd14432 : data_rom <= {16'd32195, 16'd6096};
                15'd14433 : data_rom <= {16'd32196, 16'd6093};
                15'd14434 : data_rom <= {16'd32197, 16'd6090};
                15'd14435 : data_rom <= {16'd32197, 16'd6087};
                15'd14436 : data_rom <= {16'd32198, 16'd6084};
                15'd14437 : data_rom <= {16'd32198, 16'd6081};
                15'd14438 : data_rom <= {16'd32199, 16'd6078};
                15'd14439 : data_rom <= {16'd32199, 16'd6075};
                15'd14440 : data_rom <= {16'd32200, 16'd6072};
                15'd14441 : data_rom <= {16'd32201, 16'd6068};
                15'd14442 : data_rom <= {16'd32201, 16'd6065};
                15'd14443 : data_rom <= {16'd32202, 16'd6062};
                15'd14444 : data_rom <= {16'd32202, 16'd6059};
                15'd14445 : data_rom <= {16'd32203, 16'd6056};
                15'd14446 : data_rom <= {16'd32203, 16'd6053};
                15'd14447 : data_rom <= {16'd32204, 16'd6050};
                15'd14448 : data_rom <= {16'd32205, 16'd6047};
                15'd14449 : data_rom <= {16'd32205, 16'd6044};
                15'd14450 : data_rom <= {16'd32206, 16'd6041};
                15'd14451 : data_rom <= {16'd32206, 16'd6038};
                15'd14452 : data_rom <= {16'd32207, 16'd6034};
                15'd14453 : data_rom <= {16'd32208, 16'd6031};
                15'd14454 : data_rom <= {16'd32208, 16'd6028};
                15'd14455 : data_rom <= {16'd32209, 16'd6025};
                15'd14456 : data_rom <= {16'd32209, 16'd6022};
                15'd14457 : data_rom <= {16'd32210, 16'd6019};
                15'd14458 : data_rom <= {16'd32210, 16'd6016};
                15'd14459 : data_rom <= {16'd32211, 16'd6013};
                15'd14460 : data_rom <= {16'd32212, 16'd6010};
                15'd14461 : data_rom <= {16'd32212, 16'd6007};
                15'd14462 : data_rom <= {16'd32213, 16'd6004};
                15'd14463 : data_rom <= {16'd32213, 16'd6000};
                15'd14464 : data_rom <= {16'd32214, 16'd5997};
                15'd14465 : data_rom <= {16'd32214, 16'd5994};
                15'd14466 : data_rom <= {16'd32215, 16'd5991};
                15'd14467 : data_rom <= {16'd32216, 16'd5988};
                15'd14468 : data_rom <= {16'd32216, 16'd5985};
                15'd14469 : data_rom <= {16'd32217, 16'd5982};
                15'd14470 : data_rom <= {16'd32217, 16'd5979};
                15'd14471 : data_rom <= {16'd32218, 16'd5976};
                15'd14472 : data_rom <= {16'd32218, 16'd5973};
                15'd14473 : data_rom <= {16'd32219, 16'd5970};
                15'd14474 : data_rom <= {16'd32220, 16'd5967};
                15'd14475 : data_rom <= {16'd32220, 16'd5963};
                15'd14476 : data_rom <= {16'd32221, 16'd5960};
                15'd14477 : data_rom <= {16'd32221, 16'd5957};
                15'd14478 : data_rom <= {16'd32222, 16'd5954};
                15'd14479 : data_rom <= {16'd32222, 16'd5951};
                15'd14480 : data_rom <= {16'd32223, 16'd5948};
                15'd14481 : data_rom <= {16'd32224, 16'd5945};
                15'd14482 : data_rom <= {16'd32224, 16'd5942};
                15'd14483 : data_rom <= {16'd32225, 16'd5939};
                15'd14484 : data_rom <= {16'd32225, 16'd5936};
                15'd14485 : data_rom <= {16'd32226, 16'd5933};
                15'd14486 : data_rom <= {16'd32226, 16'd5929};
                15'd14487 : data_rom <= {16'd32227, 16'd5926};
                15'd14488 : data_rom <= {16'd32228, 16'd5923};
                15'd14489 : data_rom <= {16'd32228, 16'd5920};
                15'd14490 : data_rom <= {16'd32229, 16'd5917};
                15'd14491 : data_rom <= {16'd32229, 16'd5914};
                15'd14492 : data_rom <= {16'd32230, 16'd5911};
                15'd14493 : data_rom <= {16'd32230, 16'd5908};
                15'd14494 : data_rom <= {16'd32231, 16'd5905};
                15'd14495 : data_rom <= {16'd32232, 16'd5902};
                15'd14496 : data_rom <= {16'd32232, 16'd5899};
                15'd14497 : data_rom <= {16'd32233, 16'd5895};
                15'd14498 : data_rom <= {16'd32233, 16'd5892};
                15'd14499 : data_rom <= {16'd32234, 16'd5889};
                15'd14500 : data_rom <= {16'd32234, 16'd5886};
                15'd14501 : data_rom <= {16'd32235, 16'd5883};
                15'd14502 : data_rom <= {16'd32236, 16'd5880};
                15'd14503 : data_rom <= {16'd32236, 16'd5877};
                15'd14504 : data_rom <= {16'd32237, 16'd5874};
                15'd14505 : data_rom <= {16'd32237, 16'd5871};
                15'd14506 : data_rom <= {16'd32238, 16'd5868};
                15'd14507 : data_rom <= {16'd32238, 16'd5865};
                15'd14508 : data_rom <= {16'd32239, 16'd5861};
                15'd14509 : data_rom <= {16'd32239, 16'd5858};
                15'd14510 : data_rom <= {16'd32240, 16'd5855};
                15'd14511 : data_rom <= {16'd32241, 16'd5852};
                15'd14512 : data_rom <= {16'd32241, 16'd5849};
                15'd14513 : data_rom <= {16'd32242, 16'd5846};
                15'd14514 : data_rom <= {16'd32242, 16'd5843};
                15'd14515 : data_rom <= {16'd32243, 16'd5840};
                15'd14516 : data_rom <= {16'd32243, 16'd5837};
                15'd14517 : data_rom <= {16'd32244, 16'd5834};
                15'd14518 : data_rom <= {16'd32245, 16'd5831};
                15'd14519 : data_rom <= {16'd32245, 16'd5827};
                15'd14520 : data_rom <= {16'd32246, 16'd5824};
                15'd14521 : data_rom <= {16'd32246, 16'd5821};
                15'd14522 : data_rom <= {16'd32247, 16'd5818};
                15'd14523 : data_rom <= {16'd32247, 16'd5815};
                15'd14524 : data_rom <= {16'd32248, 16'd5812};
                15'd14525 : data_rom <= {16'd32248, 16'd5809};
                15'd14526 : data_rom <= {16'd32249, 16'd5806};
                15'd14527 : data_rom <= {16'd32250, 16'd5803};
                15'd14528 : data_rom <= {16'd32250, 16'd5800};
                15'd14529 : data_rom <= {16'd32251, 16'd5797};
                15'd14530 : data_rom <= {16'd32251, 16'd5793};
                15'd14531 : data_rom <= {16'd32252, 16'd5790};
                15'd14532 : data_rom <= {16'd32252, 16'd5787};
                15'd14533 : data_rom <= {16'd32253, 16'd5784};
                15'd14534 : data_rom <= {16'd32253, 16'd5781};
                15'd14535 : data_rom <= {16'd32254, 16'd5778};
                15'd14536 : data_rom <= {16'd32255, 16'd5775};
                15'd14537 : data_rom <= {16'd32255, 16'd5772};
                15'd14538 : data_rom <= {16'd32256, 16'd5769};
                15'd14539 : data_rom <= {16'd32256, 16'd5766};
                15'd14540 : data_rom <= {16'd32257, 16'd5763};
                15'd14541 : data_rom <= {16'd32257, 16'd5759};
                15'd14542 : data_rom <= {16'd32258, 16'd5756};
                15'd14543 : data_rom <= {16'd32258, 16'd5753};
                15'd14544 : data_rom <= {16'd32259, 16'd5750};
                15'd14545 : data_rom <= {16'd32259, 16'd5747};
                15'd14546 : data_rom <= {16'd32260, 16'd5744};
                15'd14547 : data_rom <= {16'd32261, 16'd5741};
                15'd14548 : data_rom <= {16'd32261, 16'd5738};
                15'd14549 : data_rom <= {16'd32262, 16'd5735};
                15'd14550 : data_rom <= {16'd32262, 16'd5732};
                15'd14551 : data_rom <= {16'd32263, 16'd5728};
                15'd14552 : data_rom <= {16'd32263, 16'd5725};
                15'd14553 : data_rom <= {16'd32264, 16'd5722};
                15'd14554 : data_rom <= {16'd32264, 16'd5719};
                15'd14555 : data_rom <= {16'd32265, 16'd5716};
                15'd14556 : data_rom <= {16'd32266, 16'd5713};
                15'd14557 : data_rom <= {16'd32266, 16'd5710};
                15'd14558 : data_rom <= {16'd32267, 16'd5707};
                15'd14559 : data_rom <= {16'd32267, 16'd5704};
                15'd14560 : data_rom <= {16'd32268, 16'd5701};
                15'd14561 : data_rom <= {16'd32268, 16'd5698};
                15'd14562 : data_rom <= {16'd32269, 16'd5694};
                15'd14563 : data_rom <= {16'd32269, 16'd5691};
                15'd14564 : data_rom <= {16'd32270, 16'd5688};
                15'd14565 : data_rom <= {16'd32270, 16'd5685};
                15'd14566 : data_rom <= {16'd32271, 16'd5682};
                15'd14567 : data_rom <= {16'd32272, 16'd5679};
                15'd14568 : data_rom <= {16'd32272, 16'd5676};
                15'd14569 : data_rom <= {16'd32273, 16'd5673};
                15'd14570 : data_rom <= {16'd32273, 16'd5670};
                15'd14571 : data_rom <= {16'd32274, 16'd5667};
                15'd14572 : data_rom <= {16'd32274, 16'd5664};
                15'd14573 : data_rom <= {16'd32275, 16'd5660};
                15'd14574 : data_rom <= {16'd32275, 16'd5657};
                15'd14575 : data_rom <= {16'd32276, 16'd5654};
                15'd14576 : data_rom <= {16'd32276, 16'd5651};
                15'd14577 : data_rom <= {16'd32277, 16'd5648};
                15'd14578 : data_rom <= {16'd32278, 16'd5645};
                15'd14579 : data_rom <= {16'd32278, 16'd5642};
                15'd14580 : data_rom <= {16'd32279, 16'd5639};
                15'd14581 : data_rom <= {16'd32279, 16'd5636};
                15'd14582 : data_rom <= {16'd32280, 16'd5633};
                15'd14583 : data_rom <= {16'd32280, 16'd5629};
                15'd14584 : data_rom <= {16'd32281, 16'd5626};
                15'd14585 : data_rom <= {16'd32281, 16'd5623};
                15'd14586 : data_rom <= {16'd32282, 16'd5620};
                15'd14587 : data_rom <= {16'd32282, 16'd5617};
                15'd14588 : data_rom <= {16'd32283, 16'd5614};
                15'd14589 : data_rom <= {16'd32283, 16'd5611};
                15'd14590 : data_rom <= {16'd32284, 16'd5608};
                15'd14591 : data_rom <= {16'd32285, 16'd5605};
                15'd14592 : data_rom <= {16'd32285, 16'd5602};
                15'd14593 : data_rom <= {16'd32286, 16'd5599};
                15'd14594 : data_rom <= {16'd32286, 16'd5595};
                15'd14595 : data_rom <= {16'd32287, 16'd5592};
                15'd14596 : data_rom <= {16'd32287, 16'd5589};
                15'd14597 : data_rom <= {16'd32288, 16'd5586};
                15'd14598 : data_rom <= {16'd32288, 16'd5583};
                15'd14599 : data_rom <= {16'd32289, 16'd5580};
                15'd14600 : data_rom <= {16'd32289, 16'd5577};
                15'd14601 : data_rom <= {16'd32290, 16'd5574};
                15'd14602 : data_rom <= {16'd32290, 16'd5571};
                15'd14603 : data_rom <= {16'd32291, 16'd5568};
                15'd14604 : data_rom <= {16'd32291, 16'd5564};
                15'd14605 : data_rom <= {16'd32292, 16'd5561};
                15'd14606 : data_rom <= {16'd32293, 16'd5558};
                15'd14607 : data_rom <= {16'd32293, 16'd5555};
                15'd14608 : data_rom <= {16'd32294, 16'd5552};
                15'd14609 : data_rom <= {16'd32294, 16'd5549};
                15'd14610 : data_rom <= {16'd32295, 16'd5546};
                15'd14611 : data_rom <= {16'd32295, 16'd5543};
                15'd14612 : data_rom <= {16'd32296, 16'd5540};
                15'd14613 : data_rom <= {16'd32296, 16'd5537};
                15'd14614 : data_rom <= {16'd32297, 16'd5534};
                15'd14615 : data_rom <= {16'd32297, 16'd5530};
                15'd14616 : data_rom <= {16'd32298, 16'd5527};
                15'd14617 : data_rom <= {16'd32298, 16'd5524};
                15'd14618 : data_rom <= {16'd32299, 16'd5521};
                15'd14619 : data_rom <= {16'd32299, 16'd5518};
                15'd14620 : data_rom <= {16'd32300, 16'd5515};
                15'd14621 : data_rom <= {16'd32301, 16'd5512};
                15'd14622 : data_rom <= {16'd32301, 16'd5509};
                15'd14623 : data_rom <= {16'd32302, 16'd5506};
                15'd14624 : data_rom <= {16'd32302, 16'd5503};
                15'd14625 : data_rom <= {16'd32303, 16'd5499};
                15'd14626 : data_rom <= {16'd32303, 16'd5496};
                15'd14627 : data_rom <= {16'd32304, 16'd5493};
                15'd14628 : data_rom <= {16'd32304, 16'd5490};
                15'd14629 : data_rom <= {16'd32305, 16'd5487};
                15'd14630 : data_rom <= {16'd32305, 16'd5484};
                15'd14631 : data_rom <= {16'd32306, 16'd5481};
                15'd14632 : data_rom <= {16'd32306, 16'd5478};
                15'd14633 : data_rom <= {16'd32307, 16'd5475};
                15'd14634 : data_rom <= {16'd32307, 16'd5472};
                15'd14635 : data_rom <= {16'd32308, 16'd5468};
                15'd14636 : data_rom <= {16'd32308, 16'd5465};
                15'd14637 : data_rom <= {16'd32309, 16'd5462};
                15'd14638 : data_rom <= {16'd32309, 16'd5459};
                15'd14639 : data_rom <= {16'd32310, 16'd5456};
                15'd14640 : data_rom <= {16'd32311, 16'd5453};
                15'd14641 : data_rom <= {16'd32311, 16'd5450};
                15'd14642 : data_rom <= {16'd32312, 16'd5447};
                15'd14643 : data_rom <= {16'd32312, 16'd5444};
                15'd14644 : data_rom <= {16'd32313, 16'd5441};
                15'd14645 : data_rom <= {16'd32313, 16'd5437};
                15'd14646 : data_rom <= {16'd32314, 16'd5434};
                15'd14647 : data_rom <= {16'd32314, 16'd5431};
                15'd14648 : data_rom <= {16'd32315, 16'd5428};
                15'd14649 : data_rom <= {16'd32315, 16'd5425};
                15'd14650 : data_rom <= {16'd32316, 16'd5422};
                15'd14651 : data_rom <= {16'd32316, 16'd5419};
                15'd14652 : data_rom <= {16'd32317, 16'd5416};
                15'd14653 : data_rom <= {16'd32317, 16'd5413};
                15'd14654 : data_rom <= {16'd32318, 16'd5410};
                15'd14655 : data_rom <= {16'd32318, 16'd5407};
                15'd14656 : data_rom <= {16'd32319, 16'd5403};
                15'd14657 : data_rom <= {16'd32319, 16'd5400};
                15'd14658 : data_rom <= {16'd32320, 16'd5397};
                15'd14659 : data_rom <= {16'd32320, 16'd5394};
                15'd14660 : data_rom <= {16'd32321, 16'd5391};
                15'd14661 : data_rom <= {16'd32321, 16'd5388};
                15'd14662 : data_rom <= {16'd32322, 16'd5385};
                15'd14663 : data_rom <= {16'd32322, 16'd5382};
                15'd14664 : data_rom <= {16'd32323, 16'd5379};
                15'd14665 : data_rom <= {16'd32323, 16'd5376};
                15'd14666 : data_rom <= {16'd32324, 16'd5372};
                15'd14667 : data_rom <= {16'd32325, 16'd5369};
                15'd14668 : data_rom <= {16'd32325, 16'd5366};
                15'd14669 : data_rom <= {16'd32326, 16'd5363};
                15'd14670 : data_rom <= {16'd32326, 16'd5360};
                15'd14671 : data_rom <= {16'd32327, 16'd5357};
                15'd14672 : data_rom <= {16'd32327, 16'd5354};
                15'd14673 : data_rom <= {16'd32328, 16'd5351};
                15'd14674 : data_rom <= {16'd32328, 16'd5348};
                15'd14675 : data_rom <= {16'd32329, 16'd5345};
                15'd14676 : data_rom <= {16'd32329, 16'd5341};
                15'd14677 : data_rom <= {16'd32330, 16'd5338};
                15'd14678 : data_rom <= {16'd32330, 16'd5335};
                15'd14679 : data_rom <= {16'd32331, 16'd5332};
                15'd14680 : data_rom <= {16'd32331, 16'd5329};
                15'd14681 : data_rom <= {16'd32332, 16'd5326};
                15'd14682 : data_rom <= {16'd32332, 16'd5323};
                15'd14683 : data_rom <= {16'd32333, 16'd5320};
                15'd14684 : data_rom <= {16'd32333, 16'd5317};
                15'd14685 : data_rom <= {16'd32334, 16'd5314};
                15'd14686 : data_rom <= {16'd32334, 16'd5310};
                15'd14687 : data_rom <= {16'd32335, 16'd5307};
                15'd14688 : data_rom <= {16'd32335, 16'd5304};
                15'd14689 : data_rom <= {16'd32336, 16'd5301};
                15'd14690 : data_rom <= {16'd32336, 16'd5298};
                15'd14691 : data_rom <= {16'd32337, 16'd5295};
                15'd14692 : data_rom <= {16'd32337, 16'd5292};
                15'd14693 : data_rom <= {16'd32338, 16'd5289};
                15'd14694 : data_rom <= {16'd32338, 16'd5286};
                15'd14695 : data_rom <= {16'd32339, 16'd5283};
                15'd14696 : data_rom <= {16'd32339, 16'd5279};
                15'd14697 : data_rom <= {16'd32340, 16'd5276};
                15'd14698 : data_rom <= {16'd32340, 16'd5273};
                15'd14699 : data_rom <= {16'd32341, 16'd5270};
                15'd14700 : data_rom <= {16'd32341, 16'd5267};
                15'd14701 : data_rom <= {16'd32342, 16'd5264};
                15'd14702 : data_rom <= {16'd32342, 16'd5261};
                15'd14703 : data_rom <= {16'd32343, 16'd5258};
                15'd14704 : data_rom <= {16'd32343, 16'd5255};
                15'd14705 : data_rom <= {16'd32344, 16'd5252};
                15'd14706 : data_rom <= {16'd32344, 16'd5248};
                15'd14707 : data_rom <= {16'd32345, 16'd5245};
                15'd14708 : data_rom <= {16'd32345, 16'd5242};
                15'd14709 : data_rom <= {16'd32346, 16'd5239};
                15'd14710 : data_rom <= {16'd32346, 16'd5236};
                15'd14711 : data_rom <= {16'd32347, 16'd5233};
                15'd14712 : data_rom <= {16'd32347, 16'd5230};
                15'd14713 : data_rom <= {16'd32348, 16'd5227};
                15'd14714 : data_rom <= {16'd32348, 16'd5224};
                15'd14715 : data_rom <= {16'd32349, 16'd5221};
                15'd14716 : data_rom <= {16'd32349, 16'd5217};
                15'd14717 : data_rom <= {16'd32350, 16'd5214};
                15'd14718 : data_rom <= {16'd32350, 16'd5211};
                15'd14719 : data_rom <= {16'd32351, 16'd5208};
                15'd14720 : data_rom <= {16'd32351, 16'd5205};
                15'd14721 : data_rom <= {16'd32352, 16'd5202};
                15'd14722 : data_rom <= {16'd32352, 16'd5199};
                15'd14723 : data_rom <= {16'd32353, 16'd5196};
                15'd14724 : data_rom <= {16'd32353, 16'd5193};
                15'd14725 : data_rom <= {16'd32354, 16'd5189};
                15'd14726 : data_rom <= {16'd32354, 16'd5186};
                15'd14727 : data_rom <= {16'd32355, 16'd5183};
                15'd14728 : data_rom <= {16'd32355, 16'd5180};
                15'd14729 : data_rom <= {16'd32356, 16'd5177};
                15'd14730 : data_rom <= {16'd32356, 16'd5174};
                15'd14731 : data_rom <= {16'd32357, 16'd5171};
                15'd14732 : data_rom <= {16'd32357, 16'd5168};
                15'd14733 : data_rom <= {16'd32358, 16'd5165};
                15'd14734 : data_rom <= {16'd32358, 16'd5162};
                15'd14735 : data_rom <= {16'd32359, 16'd5158};
                15'd14736 : data_rom <= {16'd32359, 16'd5155};
                15'd14737 : data_rom <= {16'd32360, 16'd5152};
                15'd14738 : data_rom <= {16'd32360, 16'd5149};
                15'd14739 : data_rom <= {16'd32361, 16'd5146};
                15'd14740 : data_rom <= {16'd32361, 16'd5143};
                15'd14741 : data_rom <= {16'd32362, 16'd5140};
                15'd14742 : data_rom <= {16'd32362, 16'd5137};
                15'd14743 : data_rom <= {16'd32363, 16'd5134};
                15'd14744 : data_rom <= {16'd32363, 16'd5131};
                15'd14745 : data_rom <= {16'd32364, 16'd5127};
                15'd14746 : data_rom <= {16'd32364, 16'd5124};
                15'd14747 : data_rom <= {16'd32365, 16'd5121};
                15'd14748 : data_rom <= {16'd32365, 16'd5118};
                15'd14749 : data_rom <= {16'd32366, 16'd5115};
                15'd14750 : data_rom <= {16'd32366, 16'd5112};
                15'd14751 : data_rom <= {16'd32367, 16'd5109};
                15'd14752 : data_rom <= {16'd32367, 16'd5106};
                15'd14753 : data_rom <= {16'd32368, 16'd5103};
                15'd14754 : data_rom <= {16'd32368, 16'd5100};
                15'd14755 : data_rom <= {16'd32369, 16'd5096};
                15'd14756 : data_rom <= {16'd32369, 16'd5093};
                15'd14757 : data_rom <= {16'd32370, 16'd5090};
                15'd14758 : data_rom <= {16'd32370, 16'd5087};
                15'd14759 : data_rom <= {16'd32371, 16'd5084};
                15'd14760 : data_rom <= {16'd32371, 16'd5081};
                15'd14761 : data_rom <= {16'd32372, 16'd5078};
                15'd14762 : data_rom <= {16'd32372, 16'd5075};
                15'd14763 : data_rom <= {16'd32373, 16'd5072};
                15'd14764 : data_rom <= {16'd32373, 16'd5068};
                15'd14765 : data_rom <= {16'd32374, 16'd5065};
                15'd14766 : data_rom <= {16'd32374, 16'd5062};
                15'd14767 : data_rom <= {16'd32375, 16'd5059};
                15'd14768 : data_rom <= {16'd32375, 16'd5056};
                15'd14769 : data_rom <= {16'd32375, 16'd5053};
                15'd14770 : data_rom <= {16'd32376, 16'd5050};
                15'd14771 : data_rom <= {16'd32376, 16'd5047};
                15'd14772 : data_rom <= {16'd32377, 16'd5044};
                15'd14773 : data_rom <= {16'd32377, 16'd5041};
                15'd14774 : data_rom <= {16'd32378, 16'd5037};
                15'd14775 : data_rom <= {16'd32378, 16'd5034};
                15'd14776 : data_rom <= {16'd32379, 16'd5031};
                15'd14777 : data_rom <= {16'd32379, 16'd5028};
                15'd14778 : data_rom <= {16'd32380, 16'd5025};
                15'd14779 : data_rom <= {16'd32380, 16'd5022};
                15'd14780 : data_rom <= {16'd32381, 16'd5019};
                15'd14781 : data_rom <= {16'd32381, 16'd5016};
                15'd14782 : data_rom <= {16'd32382, 16'd5013};
                15'd14783 : data_rom <= {16'd32382, 16'd5010};
                15'd14784 : data_rom <= {16'd32383, 16'd5006};
                15'd14785 : data_rom <= {16'd32383, 16'd5003};
                15'd14786 : data_rom <= {16'd32384, 16'd5000};
                15'd14787 : data_rom <= {16'd32384, 16'd4997};
                15'd14788 : data_rom <= {16'd32385, 16'd4994};
                15'd14789 : data_rom <= {16'd32385, 16'd4991};
                15'd14790 : data_rom <= {16'd32386, 16'd4988};
                15'd14791 : data_rom <= {16'd32386, 16'd4985};
                15'd14792 : data_rom <= {16'd32387, 16'd4982};
                15'd14793 : data_rom <= {16'd32387, 16'd4978};
                15'd14794 : data_rom <= {16'd32388, 16'd4975};
                15'd14795 : data_rom <= {16'd32388, 16'd4972};
                15'd14796 : data_rom <= {16'd32388, 16'd4969};
                15'd14797 : data_rom <= {16'd32389, 16'd4966};
                15'd14798 : data_rom <= {16'd32389, 16'd4963};
                15'd14799 : data_rom <= {16'd32390, 16'd4960};
                15'd14800 : data_rom <= {16'd32390, 16'd4957};
                15'd14801 : data_rom <= {16'd32391, 16'd4954};
                15'd14802 : data_rom <= {16'd32391, 16'd4951};
                15'd14803 : data_rom <= {16'd32392, 16'd4947};
                15'd14804 : data_rom <= {16'd32392, 16'd4944};
                15'd14805 : data_rom <= {16'd32393, 16'd4941};
                15'd14806 : data_rom <= {16'd32393, 16'd4938};
                15'd14807 : data_rom <= {16'd32394, 16'd4935};
                15'd14808 : data_rom <= {16'd32394, 16'd4932};
                15'd14809 : data_rom <= {16'd32395, 16'd4929};
                15'd14810 : data_rom <= {16'd32395, 16'd4926};
                15'd14811 : data_rom <= {16'd32396, 16'd4923};
                15'd14812 : data_rom <= {16'd32396, 16'd4919};
                15'd14813 : data_rom <= {16'd32397, 16'd4916};
                15'd14814 : data_rom <= {16'd32397, 16'd4913};
                15'd14815 : data_rom <= {16'd32397, 16'd4910};
                15'd14816 : data_rom <= {16'd32398, 16'd4907};
                15'd14817 : data_rom <= {16'd32398, 16'd4904};
                15'd14818 : data_rom <= {16'd32399, 16'd4901};
                15'd14819 : data_rom <= {16'd32399, 16'd4898};
                15'd14820 : data_rom <= {16'd32400, 16'd4895};
                15'd14821 : data_rom <= {16'd32400, 16'd4891};
                15'd14822 : data_rom <= {16'd32401, 16'd4888};
                15'd14823 : data_rom <= {16'd32401, 16'd4885};
                15'd14824 : data_rom <= {16'd32402, 16'd4882};
                15'd14825 : data_rom <= {16'd32402, 16'd4879};
                15'd14826 : data_rom <= {16'd32403, 16'd4876};
                15'd14827 : data_rom <= {16'd32403, 16'd4873};
                15'd14828 : data_rom <= {16'd32404, 16'd4870};
                15'd14829 : data_rom <= {16'd32404, 16'd4867};
                15'd14830 : data_rom <= {16'd32404, 16'd4864};
                15'd14831 : data_rom <= {16'd32405, 16'd4860};
                15'd14832 : data_rom <= {16'd32405, 16'd4857};
                15'd14833 : data_rom <= {16'd32406, 16'd4854};
                15'd14834 : data_rom <= {16'd32406, 16'd4851};
                15'd14835 : data_rom <= {16'd32407, 16'd4848};
                15'd14836 : data_rom <= {16'd32407, 16'd4845};
                15'd14837 : data_rom <= {16'd32408, 16'd4842};
                15'd14838 : data_rom <= {16'd32408, 16'd4839};
                15'd14839 : data_rom <= {16'd32409, 16'd4836};
                15'd14840 : data_rom <= {16'd32409, 16'd4832};
                15'd14841 : data_rom <= {16'd32410, 16'd4829};
                15'd14842 : data_rom <= {16'd32410, 16'd4826};
                15'd14843 : data_rom <= {16'd32411, 16'd4823};
                15'd14844 : data_rom <= {16'd32411, 16'd4820};
                15'd14845 : data_rom <= {16'd32411, 16'd4817};
                15'd14846 : data_rom <= {16'd32412, 16'd4814};
                15'd14847 : data_rom <= {16'd32412, 16'd4811};
                15'd14848 : data_rom <= {16'd32413, 16'd4808};
                15'd14849 : data_rom <= {16'd32413, 16'd4805};
                15'd14850 : data_rom <= {16'd32414, 16'd4801};
                15'd14851 : data_rom <= {16'd32414, 16'd4798};
                15'd14852 : data_rom <= {16'd32415, 16'd4795};
                15'd14853 : data_rom <= {16'd32415, 16'd4792};
                15'd14854 : data_rom <= {16'd32416, 16'd4789};
                15'd14855 : data_rom <= {16'd32416, 16'd4786};
                15'd14856 : data_rom <= {16'd32417, 16'd4783};
                15'd14857 : data_rom <= {16'd32417, 16'd4780};
                15'd14858 : data_rom <= {16'd32417, 16'd4777};
                15'd14859 : data_rom <= {16'd32418, 16'd4773};
                15'd14860 : data_rom <= {16'd32418, 16'd4770};
                15'd14861 : data_rom <= {16'd32419, 16'd4767};
                15'd14862 : data_rom <= {16'd32419, 16'd4764};
                15'd14863 : data_rom <= {16'd32420, 16'd4761};
                15'd14864 : data_rom <= {16'd32420, 16'd4758};
                15'd14865 : data_rom <= {16'd32421, 16'd4755};
                15'd14866 : data_rom <= {16'd32421, 16'd4752};
                15'd14867 : data_rom <= {16'd32422, 16'd4749};
                15'd14868 : data_rom <= {16'd32422, 16'd4745};
                15'd14869 : data_rom <= {16'd32422, 16'd4742};
                15'd14870 : data_rom <= {16'd32423, 16'd4739};
                15'd14871 : data_rom <= {16'd32423, 16'd4736};
                15'd14872 : data_rom <= {16'd32424, 16'd4733};
                15'd14873 : data_rom <= {16'd32424, 16'd4730};
                15'd14874 : data_rom <= {16'd32425, 16'd4727};
                15'd14875 : data_rom <= {16'd32425, 16'd4724};
                15'd14876 : data_rom <= {16'd32426, 16'd4721};
                15'd14877 : data_rom <= {16'd32426, 16'd4717};
                15'd14878 : data_rom <= {16'd32427, 16'd4714};
                15'd14879 : data_rom <= {16'd32427, 16'd4711};
                15'd14880 : data_rom <= {16'd32427, 16'd4708};
                15'd14881 : data_rom <= {16'd32428, 16'd4705};
                15'd14882 : data_rom <= {16'd32428, 16'd4702};
                15'd14883 : data_rom <= {16'd32429, 16'd4699};
                15'd14884 : data_rom <= {16'd32429, 16'd4696};
                15'd14885 : data_rom <= {16'd32430, 16'd4693};
                15'd14886 : data_rom <= {16'd32430, 16'd4689};
                15'd14887 : data_rom <= {16'd32431, 16'd4686};
                15'd14888 : data_rom <= {16'd32431, 16'd4683};
                15'd14889 : data_rom <= {16'd32431, 16'd4680};
                15'd14890 : data_rom <= {16'd32432, 16'd4677};
                15'd14891 : data_rom <= {16'd32432, 16'd4674};
                15'd14892 : data_rom <= {16'd32433, 16'd4671};
                15'd14893 : data_rom <= {16'd32433, 16'd4668};
                15'd14894 : data_rom <= {16'd32434, 16'd4665};
                15'd14895 : data_rom <= {16'd32434, 16'd4662};
                15'd14896 : data_rom <= {16'd32435, 16'd4658};
                15'd14897 : data_rom <= {16'd32435, 16'd4655};
                15'd14898 : data_rom <= {16'd32436, 16'd4652};
                15'd14899 : data_rom <= {16'd32436, 16'd4649};
                15'd14900 : data_rom <= {16'd32436, 16'd4646};
                15'd14901 : data_rom <= {16'd32437, 16'd4643};
                15'd14902 : data_rom <= {16'd32437, 16'd4640};
                15'd14903 : data_rom <= {16'd32438, 16'd4637};
                15'd14904 : data_rom <= {16'd32438, 16'd4634};
                15'd14905 : data_rom <= {16'd32439, 16'd4630};
                15'd14906 : data_rom <= {16'd32439, 16'd4627};
                15'd14907 : data_rom <= {16'd32440, 16'd4624};
                15'd14908 : data_rom <= {16'd32440, 16'd4621};
                15'd14909 : data_rom <= {16'd32440, 16'd4618};
                15'd14910 : data_rom <= {16'd32441, 16'd4615};
                15'd14911 : data_rom <= {16'd32441, 16'd4612};
                15'd14912 : data_rom <= {16'd32442, 16'd4609};
                15'd14913 : data_rom <= {16'd32442, 16'd4606};
                15'd14914 : data_rom <= {16'd32443, 16'd4602};
                15'd14915 : data_rom <= {16'd32443, 16'd4599};
                15'd14916 : data_rom <= {16'd32443, 16'd4596};
                15'd14917 : data_rom <= {16'd32444, 16'd4593};
                15'd14918 : data_rom <= {16'd32444, 16'd4590};
                15'd14919 : data_rom <= {16'd32445, 16'd4587};
                15'd14920 : data_rom <= {16'd32445, 16'd4584};
                15'd14921 : data_rom <= {16'd32446, 16'd4581};
                15'd14922 : data_rom <= {16'd32446, 16'd4578};
                15'd14923 : data_rom <= {16'd32447, 16'd4574};
                15'd14924 : data_rom <= {16'd32447, 16'd4571};
                15'd14925 : data_rom <= {16'd32447, 16'd4568};
                15'd14926 : data_rom <= {16'd32448, 16'd4565};
                15'd14927 : data_rom <= {16'd32448, 16'd4562};
                15'd14928 : data_rom <= {16'd32449, 16'd4559};
                15'd14929 : data_rom <= {16'd32449, 16'd4556};
                15'd14930 : data_rom <= {16'd32450, 16'd4553};
                15'd14931 : data_rom <= {16'd32450, 16'd4550};
                15'd14932 : data_rom <= {16'd32450, 16'd4546};
                15'd14933 : data_rom <= {16'd32451, 16'd4543};
                15'd14934 : data_rom <= {16'd32451, 16'd4540};
                15'd14935 : data_rom <= {16'd32452, 16'd4537};
                15'd14936 : data_rom <= {16'd32452, 16'd4534};
                15'd14937 : data_rom <= {16'd32453, 16'd4531};
                15'd14938 : data_rom <= {16'd32453, 16'd4528};
                15'd14939 : data_rom <= {16'd32454, 16'd4525};
                15'd14940 : data_rom <= {16'd32454, 16'd4522};
                15'd14941 : data_rom <= {16'd32454, 16'd4518};
                15'd14942 : data_rom <= {16'd32455, 16'd4515};
                15'd14943 : data_rom <= {16'd32455, 16'd4512};
                15'd14944 : data_rom <= {16'd32456, 16'd4509};
                15'd14945 : data_rom <= {16'd32456, 16'd4506};
                15'd14946 : data_rom <= {16'd32457, 16'd4503};
                15'd14947 : data_rom <= {16'd32457, 16'd4500};
                15'd14948 : data_rom <= {16'd32457, 16'd4497};
                15'd14949 : data_rom <= {16'd32458, 16'd4494};
                15'd14950 : data_rom <= {16'd32458, 16'd4490};
                15'd14951 : data_rom <= {16'd32459, 16'd4487};
                15'd14952 : data_rom <= {16'd32459, 16'd4484};
                15'd14953 : data_rom <= {16'd32460, 16'd4481};
                15'd14954 : data_rom <= {16'd32460, 16'd4478};
                15'd14955 : data_rom <= {16'd32460, 16'd4475};
                15'd14956 : data_rom <= {16'd32461, 16'd4472};
                15'd14957 : data_rom <= {16'd32461, 16'd4469};
                15'd14958 : data_rom <= {16'd32462, 16'd4466};
                15'd14959 : data_rom <= {16'd32462, 16'd4462};
                15'd14960 : data_rom <= {16'd32463, 16'd4459};
                15'd14961 : data_rom <= {16'd32463, 16'd4456};
                15'd14962 : data_rom <= {16'd32463, 16'd4453};
                15'd14963 : data_rom <= {16'd32464, 16'd4450};
                15'd14964 : data_rom <= {16'd32464, 16'd4447};
                15'd14965 : data_rom <= {16'd32465, 16'd4444};
                15'd14966 : data_rom <= {16'd32465, 16'd4441};
                15'd14967 : data_rom <= {16'd32466, 16'd4438};
                15'd14968 : data_rom <= {16'd32466, 16'd4434};
                15'd14969 : data_rom <= {16'd32466, 16'd4431};
                15'd14970 : data_rom <= {16'd32467, 16'd4428};
                15'd14971 : data_rom <= {16'd32467, 16'd4425};
                15'd14972 : data_rom <= {16'd32468, 16'd4422};
                15'd14973 : data_rom <= {16'd32468, 16'd4419};
                15'd14974 : data_rom <= {16'd32469, 16'd4416};
                15'd14975 : data_rom <= {16'd32469, 16'd4413};
                15'd14976 : data_rom <= {16'd32469, 16'd4409};
                15'd14977 : data_rom <= {16'd32470, 16'd4406};
                15'd14978 : data_rom <= {16'd32470, 16'd4403};
                15'd14979 : data_rom <= {16'd32471, 16'd4400};
                15'd14980 : data_rom <= {16'd32471, 16'd4397};
                15'd14981 : data_rom <= {16'd32472, 16'd4394};
                15'd14982 : data_rom <= {16'd32472, 16'd4391};
                15'd14983 : data_rom <= {16'd32472, 16'd4388};
                15'd14984 : data_rom <= {16'd32473, 16'd4385};
                15'd14985 : data_rom <= {16'd32473, 16'd4381};
                15'd14986 : data_rom <= {16'd32474, 16'd4378};
                15'd14987 : data_rom <= {16'd32474, 16'd4375};
                15'd14988 : data_rom <= {16'd32474, 16'd4372};
                15'd14989 : data_rom <= {16'd32475, 16'd4369};
                15'd14990 : data_rom <= {16'd32475, 16'd4366};
                15'd14991 : data_rom <= {16'd32476, 16'd4363};
                15'd14992 : data_rom <= {16'd32476, 16'd4360};
                15'd14993 : data_rom <= {16'd32477, 16'd4357};
                15'd14994 : data_rom <= {16'd32477, 16'd4353};
                15'd14995 : data_rom <= {16'd32477, 16'd4350};
                15'd14996 : data_rom <= {16'd32478, 16'd4347};
                15'd14997 : data_rom <= {16'd32478, 16'd4344};
                15'd14998 : data_rom <= {16'd32479, 16'd4341};
                15'd14999 : data_rom <= {16'd32479, 16'd4338};
                15'd15000 : data_rom <= {16'd32479, 16'd4335};
                15'd15001 : data_rom <= {16'd32480, 16'd4332};
                15'd15002 : data_rom <= {16'd32480, 16'd4329};
                15'd15003 : data_rom <= {16'd32481, 16'd4325};
                15'd15004 : data_rom <= {16'd32481, 16'd4322};
                15'd15005 : data_rom <= {16'd32482, 16'd4319};
                15'd15006 : data_rom <= {16'd32482, 16'd4316};
                15'd15007 : data_rom <= {16'd32482, 16'd4313};
                15'd15008 : data_rom <= {16'd32483, 16'd4310};
                15'd15009 : data_rom <= {16'd32483, 16'd4307};
                15'd15010 : data_rom <= {16'd32484, 16'd4304};
                15'd15011 : data_rom <= {16'd32484, 16'd4301};
                15'd15012 : data_rom <= {16'd32484, 16'd4297};
                15'd15013 : data_rom <= {16'd32485, 16'd4294};
                15'd15014 : data_rom <= {16'd32485, 16'd4291};
                15'd15015 : data_rom <= {16'd32486, 16'd4288};
                15'd15016 : data_rom <= {16'd32486, 16'd4285};
                15'd15017 : data_rom <= {16'd32486, 16'd4282};
                15'd15018 : data_rom <= {16'd32487, 16'd4279};
                15'd15019 : data_rom <= {16'd32487, 16'd4276};
                15'd15020 : data_rom <= {16'd32488, 16'd4272};
                15'd15021 : data_rom <= {16'd32488, 16'd4269};
                15'd15022 : data_rom <= {16'd32489, 16'd4266};
                15'd15023 : data_rom <= {16'd32489, 16'd4263};
                15'd15024 : data_rom <= {16'd32489, 16'd4260};
                15'd15025 : data_rom <= {16'd32490, 16'd4257};
                15'd15026 : data_rom <= {16'd32490, 16'd4254};
                15'd15027 : data_rom <= {16'd32491, 16'd4251};
                15'd15028 : data_rom <= {16'd32491, 16'd4248};
                15'd15029 : data_rom <= {16'd32491, 16'd4244};
                15'd15030 : data_rom <= {16'd32492, 16'd4241};
                15'd15031 : data_rom <= {16'd32492, 16'd4238};
                15'd15032 : data_rom <= {16'd32493, 16'd4235};
                15'd15033 : data_rom <= {16'd32493, 16'd4232};
                15'd15034 : data_rom <= {16'd32493, 16'd4229};
                15'd15035 : data_rom <= {16'd32494, 16'd4226};
                15'd15036 : data_rom <= {16'd32494, 16'd4223};
                15'd15037 : data_rom <= {16'd32495, 16'd4220};
                15'd15038 : data_rom <= {16'd32495, 16'd4216};
                15'd15039 : data_rom <= {16'd32495, 16'd4213};
                15'd15040 : data_rom <= {16'd32496, 16'd4210};
                15'd15041 : data_rom <= {16'd32496, 16'd4207};
                15'd15042 : data_rom <= {16'd32497, 16'd4204};
                15'd15043 : data_rom <= {16'd32497, 16'd4201};
                15'd15044 : data_rom <= {16'd32497, 16'd4198};
                15'd15045 : data_rom <= {16'd32498, 16'd4195};
                15'd15046 : data_rom <= {16'd32498, 16'd4191};
                15'd15047 : data_rom <= {16'd32499, 16'd4188};
                15'd15048 : data_rom <= {16'd32499, 16'd4185};
                15'd15049 : data_rom <= {16'd32499, 16'd4182};
                15'd15050 : data_rom <= {16'd32500, 16'd4179};
                15'd15051 : data_rom <= {16'd32500, 16'd4176};
                15'd15052 : data_rom <= {16'd32501, 16'd4173};
                15'd15053 : data_rom <= {16'd32501, 16'd4170};
                15'd15054 : data_rom <= {16'd32501, 16'd4167};
                15'd15055 : data_rom <= {16'd32502, 16'd4163};
                15'd15056 : data_rom <= {16'd32502, 16'd4160};
                15'd15057 : data_rom <= {16'd32503, 16'd4157};
                15'd15058 : data_rom <= {16'd32503, 16'd4154};
                15'd15059 : data_rom <= {16'd32503, 16'd4151};
                15'd15060 : data_rom <= {16'd32504, 16'd4148};
                15'd15061 : data_rom <= {16'd32504, 16'd4145};
                15'd15062 : data_rom <= {16'd32505, 16'd4142};
                15'd15063 : data_rom <= {16'd32505, 16'd4139};
                15'd15064 : data_rom <= {16'd32505, 16'd4135};
                15'd15065 : data_rom <= {16'd32506, 16'd4132};
                15'd15066 : data_rom <= {16'd32506, 16'd4129};
                15'd15067 : data_rom <= {16'd32507, 16'd4126};
                15'd15068 : data_rom <= {16'd32507, 16'd4123};
                15'd15069 : data_rom <= {16'd32507, 16'd4120};
                15'd15070 : data_rom <= {16'd32508, 16'd4117};
                15'd15071 : data_rom <= {16'd32508, 16'd4114};
                15'd15072 : data_rom <= {16'd32509, 16'd4110};
                15'd15073 : data_rom <= {16'd32509, 16'd4107};
                15'd15074 : data_rom <= {16'd32509, 16'd4104};
                15'd15075 : data_rom <= {16'd32510, 16'd4101};
                15'd15076 : data_rom <= {16'd32510, 16'd4098};
                15'd15077 : data_rom <= {16'd32511, 16'd4095};
                15'd15078 : data_rom <= {16'd32511, 16'd4092};
                15'd15079 : data_rom <= {16'd32511, 16'd4089};
                15'd15080 : data_rom <= {16'd32512, 16'd4086};
                15'd15081 : data_rom <= {16'd32512, 16'd4082};
                15'd15082 : data_rom <= {16'd32513, 16'd4079};
                15'd15083 : data_rom <= {16'd32513, 16'd4076};
                15'd15084 : data_rom <= {16'd32513, 16'd4073};
                15'd15085 : data_rom <= {16'd32514, 16'd4070};
                15'd15086 : data_rom <= {16'd32514, 16'd4067};
                15'd15087 : data_rom <= {16'd32514, 16'd4064};
                15'd15088 : data_rom <= {16'd32515, 16'd4061};
                15'd15089 : data_rom <= {16'd32515, 16'd4057};
                15'd15090 : data_rom <= {16'd32516, 16'd4054};
                15'd15091 : data_rom <= {16'd32516, 16'd4051};
                15'd15092 : data_rom <= {16'd32516, 16'd4048};
                15'd15093 : data_rom <= {16'd32517, 16'd4045};
                15'd15094 : data_rom <= {16'd32517, 16'd4042};
                15'd15095 : data_rom <= {16'd32518, 16'd4039};
                15'd15096 : data_rom <= {16'd32518, 16'd4036};
                15'd15097 : data_rom <= {16'd32518, 16'd4033};
                15'd15098 : data_rom <= {16'd32519, 16'd4029};
                15'd15099 : data_rom <= {16'd32519, 16'd4026};
                15'd15100 : data_rom <= {16'd32520, 16'd4023};
                15'd15101 : data_rom <= {16'd32520, 16'd4020};
                15'd15102 : data_rom <= {16'd32520, 16'd4017};
                15'd15103 : data_rom <= {16'd32521, 16'd4014};
                15'd15104 : data_rom <= {16'd32521, 16'd4011};
                15'd15105 : data_rom <= {16'd32521, 16'd4008};
                15'd15106 : data_rom <= {16'd32522, 16'd4004};
                15'd15107 : data_rom <= {16'd32522, 16'd4001};
                15'd15108 : data_rom <= {16'd32523, 16'd3998};
                15'd15109 : data_rom <= {16'd32523, 16'd3995};
                15'd15110 : data_rom <= {16'd32523, 16'd3992};
                15'd15111 : data_rom <= {16'd32524, 16'd3989};
                15'd15112 : data_rom <= {16'd32524, 16'd3986};
                15'd15113 : data_rom <= {16'd32525, 16'd3983};
                15'd15114 : data_rom <= {16'd32525, 16'd3980};
                15'd15115 : data_rom <= {16'd32525, 16'd3976};
                15'd15116 : data_rom <= {16'd32526, 16'd3973};
                15'd15117 : data_rom <= {16'd32526, 16'd3970};
                15'd15118 : data_rom <= {16'd32526, 16'd3967};
                15'd15119 : data_rom <= {16'd32527, 16'd3964};
                15'd15120 : data_rom <= {16'd32527, 16'd3961};
                15'd15121 : data_rom <= {16'd32528, 16'd3958};
                15'd15122 : data_rom <= {16'd32528, 16'd3955};
                15'd15123 : data_rom <= {16'd32528, 16'd3951};
                15'd15124 : data_rom <= {16'd32529, 16'd3948};
                15'd15125 : data_rom <= {16'd32529, 16'd3945};
                15'd15126 : data_rom <= {16'd32529, 16'd3942};
                15'd15127 : data_rom <= {16'd32530, 16'd3939};
                15'd15128 : data_rom <= {16'd32530, 16'd3936};
                15'd15129 : data_rom <= {16'd32531, 16'd3933};
                15'd15130 : data_rom <= {16'd32531, 16'd3930};
                15'd15131 : data_rom <= {16'd32531, 16'd3926};
                15'd15132 : data_rom <= {16'd32532, 16'd3923};
                15'd15133 : data_rom <= {16'd32532, 16'd3920};
                15'd15134 : data_rom <= {16'd32532, 16'd3917};
                15'd15135 : data_rom <= {16'd32533, 16'd3914};
                15'd15136 : data_rom <= {16'd32533, 16'd3911};
                15'd15137 : data_rom <= {16'd32534, 16'd3908};
                15'd15138 : data_rom <= {16'd32534, 16'd3905};
                15'd15139 : data_rom <= {16'd32534, 16'd3902};
                15'd15140 : data_rom <= {16'd32535, 16'd3898};
                15'd15141 : data_rom <= {16'd32535, 16'd3895};
                15'd15142 : data_rom <= {16'd32535, 16'd3892};
                15'd15143 : data_rom <= {16'd32536, 16'd3889};
                15'd15144 : data_rom <= {16'd32536, 16'd3886};
                15'd15145 : data_rom <= {16'd32537, 16'd3883};
                15'd15146 : data_rom <= {16'd32537, 16'd3880};
                15'd15147 : data_rom <= {16'd32537, 16'd3877};
                15'd15148 : data_rom <= {16'd32538, 16'd3873};
                15'd15149 : data_rom <= {16'd32538, 16'd3870};
                15'd15150 : data_rom <= {16'd32538, 16'd3867};
                15'd15151 : data_rom <= {16'd32539, 16'd3864};
                15'd15152 : data_rom <= {16'd32539, 16'd3861};
                15'd15153 : data_rom <= {16'd32540, 16'd3858};
                15'd15154 : data_rom <= {16'd32540, 16'd3855};
                15'd15155 : data_rom <= {16'd32540, 16'd3852};
                15'd15156 : data_rom <= {16'd32541, 16'd3849};
                15'd15157 : data_rom <= {16'd32541, 16'd3845};
                15'd15158 : data_rom <= {16'd32541, 16'd3842};
                15'd15159 : data_rom <= {16'd32542, 16'd3839};
                15'd15160 : data_rom <= {16'd32542, 16'd3836};
                15'd15161 : data_rom <= {16'd32542, 16'd3833};
                15'd15162 : data_rom <= {16'd32543, 16'd3830};
                15'd15163 : data_rom <= {16'd32543, 16'd3827};
                15'd15164 : data_rom <= {16'd32544, 16'd3824};
                15'd15165 : data_rom <= {16'd32544, 16'd3820};
                15'd15166 : data_rom <= {16'd32544, 16'd3817};
                15'd15167 : data_rom <= {16'd32545, 16'd3814};
                15'd15168 : data_rom <= {16'd32545, 16'd3811};
                15'd15169 : data_rom <= {16'd32545, 16'd3808};
                15'd15170 : data_rom <= {16'd32546, 16'd3805};
                15'd15171 : data_rom <= {16'd32546, 16'd3802};
                15'd15172 : data_rom <= {16'd32547, 16'd3799};
                15'd15173 : data_rom <= {16'd32547, 16'd3795};
                15'd15174 : data_rom <= {16'd32547, 16'd3792};
                15'd15175 : data_rom <= {16'd32548, 16'd3789};
                15'd15176 : data_rom <= {16'd32548, 16'd3786};
                15'd15177 : data_rom <= {16'd32548, 16'd3783};
                15'd15178 : data_rom <= {16'd32549, 16'd3780};
                15'd15179 : data_rom <= {16'd32549, 16'd3777};
                15'd15180 : data_rom <= {16'd32549, 16'd3774};
                15'd15181 : data_rom <= {16'd32550, 16'd3771};
                15'd15182 : data_rom <= {16'd32550, 16'd3767};
                15'd15183 : data_rom <= {16'd32551, 16'd3764};
                15'd15184 : data_rom <= {16'd32551, 16'd3761};
                15'd15185 : data_rom <= {16'd32551, 16'd3758};
                15'd15186 : data_rom <= {16'd32552, 16'd3755};
                15'd15187 : data_rom <= {16'd32552, 16'd3752};
                15'd15188 : data_rom <= {16'd32552, 16'd3749};
                15'd15189 : data_rom <= {16'd32553, 16'd3746};
                15'd15190 : data_rom <= {16'd32553, 16'd3742};
                15'd15191 : data_rom <= {16'd32553, 16'd3739};
                15'd15192 : data_rom <= {16'd32554, 16'd3736};
                15'd15193 : data_rom <= {16'd32554, 16'd3733};
                15'd15194 : data_rom <= {16'd32554, 16'd3730};
                15'd15195 : data_rom <= {16'd32555, 16'd3727};
                15'd15196 : data_rom <= {16'd32555, 16'd3724};
                15'd15197 : data_rom <= {16'd32556, 16'd3721};
                15'd15198 : data_rom <= {16'd32556, 16'd3717};
                15'd15199 : data_rom <= {16'd32556, 16'd3714};
                15'd15200 : data_rom <= {16'd32557, 16'd3711};
                15'd15201 : data_rom <= {16'd32557, 16'd3708};
                15'd15202 : data_rom <= {16'd32557, 16'd3705};
                15'd15203 : data_rom <= {16'd32558, 16'd3702};
                15'd15204 : data_rom <= {16'd32558, 16'd3699};
                15'd15205 : data_rom <= {16'd32558, 16'd3696};
                15'd15206 : data_rom <= {16'd32559, 16'd3692};
                15'd15207 : data_rom <= {16'd32559, 16'd3689};
                15'd15208 : data_rom <= {16'd32559, 16'd3686};
                15'd15209 : data_rom <= {16'd32560, 16'd3683};
                15'd15210 : data_rom <= {16'd32560, 16'd3680};
                15'd15211 : data_rom <= {16'd32561, 16'd3677};
                15'd15212 : data_rom <= {16'd32561, 16'd3674};
                15'd15213 : data_rom <= {16'd32561, 16'd3671};
                15'd15214 : data_rom <= {16'd32562, 16'd3668};
                15'd15215 : data_rom <= {16'd32562, 16'd3664};
                15'd15216 : data_rom <= {16'd32562, 16'd3661};
                15'd15217 : data_rom <= {16'd32563, 16'd3658};
                15'd15218 : data_rom <= {16'd32563, 16'd3655};
                15'd15219 : data_rom <= {16'd32563, 16'd3652};
                15'd15220 : data_rom <= {16'd32564, 16'd3649};
                15'd15221 : data_rom <= {16'd32564, 16'd3646};
                15'd15222 : data_rom <= {16'd32564, 16'd3643};
                15'd15223 : data_rom <= {16'd32565, 16'd3639};
                15'd15224 : data_rom <= {16'd32565, 16'd3636};
                15'd15225 : data_rom <= {16'd32565, 16'd3633};
                15'd15226 : data_rom <= {16'd32566, 16'd3630};
                15'd15227 : data_rom <= {16'd32566, 16'd3627};
                15'd15228 : data_rom <= {16'd32566, 16'd3624};
                15'd15229 : data_rom <= {16'd32567, 16'd3621};
                15'd15230 : data_rom <= {16'd32567, 16'd3618};
                15'd15231 : data_rom <= {16'd32567, 16'd3614};
                15'd15232 : data_rom <= {16'd32568, 16'd3611};
                15'd15233 : data_rom <= {16'd32568, 16'd3608};
                15'd15234 : data_rom <= {16'd32569, 16'd3605};
                15'd15235 : data_rom <= {16'd32569, 16'd3602};
                15'd15236 : data_rom <= {16'd32569, 16'd3599};
                15'd15237 : data_rom <= {16'd32570, 16'd3596};
                15'd15238 : data_rom <= {16'd32570, 16'd3593};
                15'd15239 : data_rom <= {16'd32570, 16'd3589};
                15'd15240 : data_rom <= {16'd32571, 16'd3586};
                15'd15241 : data_rom <= {16'd32571, 16'd3583};
                15'd15242 : data_rom <= {16'd32571, 16'd3580};
                15'd15243 : data_rom <= {16'd32572, 16'd3577};
                15'd15244 : data_rom <= {16'd32572, 16'd3574};
                15'd15245 : data_rom <= {16'd32572, 16'd3571};
                15'd15246 : data_rom <= {16'd32573, 16'd3568};
                15'd15247 : data_rom <= {16'd32573, 16'd3564};
                15'd15248 : data_rom <= {16'd32573, 16'd3561};
                15'd15249 : data_rom <= {16'd32574, 16'd3558};
                15'd15250 : data_rom <= {16'd32574, 16'd3555};
                15'd15251 : data_rom <= {16'd32574, 16'd3552};
                15'd15252 : data_rom <= {16'd32575, 16'd3549};
                15'd15253 : data_rom <= {16'd32575, 16'd3546};
                15'd15254 : data_rom <= {16'd32575, 16'd3543};
                15'd15255 : data_rom <= {16'd32576, 16'd3539};
                15'd15256 : data_rom <= {16'd32576, 16'd3536};
                15'd15257 : data_rom <= {16'd32576, 16'd3533};
                15'd15258 : data_rom <= {16'd32577, 16'd3530};
                15'd15259 : data_rom <= {16'd32577, 16'd3527};
                15'd15260 : data_rom <= {16'd32577, 16'd3524};
                15'd15261 : data_rom <= {16'd32578, 16'd3521};
                15'd15262 : data_rom <= {16'd32578, 16'd3518};
                15'd15263 : data_rom <= {16'd32578, 16'd3514};
                15'd15264 : data_rom <= {16'd32579, 16'd3511};
                15'd15265 : data_rom <= {16'd32579, 16'd3508};
                15'd15266 : data_rom <= {16'd32579, 16'd3505};
                15'd15267 : data_rom <= {16'd32580, 16'd3502};
                15'd15268 : data_rom <= {16'd32580, 16'd3499};
                15'd15269 : data_rom <= {16'd32580, 16'd3496};
                15'd15270 : data_rom <= {16'd32581, 16'd3493};
                15'd15271 : data_rom <= {16'd32581, 16'd3490};
                15'd15272 : data_rom <= {16'd32581, 16'd3486};
                15'd15273 : data_rom <= {16'd32582, 16'd3483};
                15'd15274 : data_rom <= {16'd32582, 16'd3480};
                15'd15275 : data_rom <= {16'd32582, 16'd3477};
                15'd15276 : data_rom <= {16'd32583, 16'd3474};
                15'd15277 : data_rom <= {16'd32583, 16'd3471};
                15'd15278 : data_rom <= {16'd32583, 16'd3468};
                15'd15279 : data_rom <= {16'd32584, 16'd3465};
                15'd15280 : data_rom <= {16'd32584, 16'd3461};
                15'd15281 : data_rom <= {16'd32584, 16'd3458};
                15'd15282 : data_rom <= {16'd32585, 16'd3455};
                15'd15283 : data_rom <= {16'd32585, 16'd3452};
                15'd15284 : data_rom <= {16'd32585, 16'd3449};
                15'd15285 : data_rom <= {16'd32586, 16'd3446};
                15'd15286 : data_rom <= {16'd32586, 16'd3443};
                15'd15287 : data_rom <= {16'd32586, 16'd3440};
                15'd15288 : data_rom <= {16'd32587, 16'd3436};
                15'd15289 : data_rom <= {16'd32587, 16'd3433};
                15'd15290 : data_rom <= {16'd32587, 16'd3430};
                15'd15291 : data_rom <= {16'd32588, 16'd3427};
                15'd15292 : data_rom <= {16'd32588, 16'd3424};
                15'd15293 : data_rom <= {16'd32588, 16'd3421};
                15'd15294 : data_rom <= {16'd32589, 16'd3418};
                15'd15295 : data_rom <= {16'd32589, 16'd3415};
                15'd15296 : data_rom <= {16'd32589, 16'd3411};
                15'd15297 : data_rom <= {16'd32590, 16'd3408};
                15'd15298 : data_rom <= {16'd32590, 16'd3405};
                15'd15299 : data_rom <= {16'd32590, 16'd3402};
                15'd15300 : data_rom <= {16'd32591, 16'd3399};
                15'd15301 : data_rom <= {16'd32591, 16'd3396};
                15'd15302 : data_rom <= {16'd32591, 16'd3393};
                15'd15303 : data_rom <= {16'd32592, 16'd3390};
                15'd15304 : data_rom <= {16'd32592, 16'd3386};
                15'd15305 : data_rom <= {16'd32592, 16'd3383};
                15'd15306 : data_rom <= {16'd32593, 16'd3380};
                15'd15307 : data_rom <= {16'd32593, 16'd3377};
                15'd15308 : data_rom <= {16'd32593, 16'd3374};
                15'd15309 : data_rom <= {16'd32594, 16'd3371};
                15'd15310 : data_rom <= {16'd32594, 16'd3368};
                15'd15311 : data_rom <= {16'd32594, 16'd3365};
                15'd15312 : data_rom <= {16'd32595, 16'd3361};
                15'd15313 : data_rom <= {16'd32595, 16'd3358};
                15'd15314 : data_rom <= {16'd32595, 16'd3355};
                15'd15315 : data_rom <= {16'd32596, 16'd3352};
                15'd15316 : data_rom <= {16'd32596, 16'd3349};
                15'd15317 : data_rom <= {16'd32596, 16'd3346};
                15'd15318 : data_rom <= {16'd32597, 16'd3343};
                15'd15319 : data_rom <= {16'd32597, 16'd3340};
                15'd15320 : data_rom <= {16'd32597, 16'd3336};
                15'd15321 : data_rom <= {16'd32597, 16'd3333};
                15'd15322 : data_rom <= {16'd32598, 16'd3330};
                15'd15323 : data_rom <= {16'd32598, 16'd3327};
                15'd15324 : data_rom <= {16'd32598, 16'd3324};
                15'd15325 : data_rom <= {16'd32599, 16'd3321};
                15'd15326 : data_rom <= {16'd32599, 16'd3318};
                15'd15327 : data_rom <= {16'd32599, 16'd3315};
                15'd15328 : data_rom <= {16'd32600, 16'd3311};
                15'd15329 : data_rom <= {16'd32600, 16'd3308};
                15'd15330 : data_rom <= {16'd32600, 16'd3305};
                15'd15331 : data_rom <= {16'd32601, 16'd3302};
                15'd15332 : data_rom <= {16'd32601, 16'd3299};
                15'd15333 : data_rom <= {16'd32601, 16'd3296};
                15'd15334 : data_rom <= {16'd32602, 16'd3293};
                15'd15335 : data_rom <= {16'd32602, 16'd3290};
                15'd15336 : data_rom <= {16'd32602, 16'd3286};
                15'd15337 : data_rom <= {16'd32603, 16'd3283};
                15'd15338 : data_rom <= {16'd32603, 16'd3280};
                15'd15339 : data_rom <= {16'd32603, 16'd3277};
                15'd15340 : data_rom <= {16'd32603, 16'd3274};
                15'd15341 : data_rom <= {16'd32604, 16'd3271};
                15'd15342 : data_rom <= {16'd32604, 16'd3268};
                15'd15343 : data_rom <= {16'd32604, 16'd3265};
                15'd15344 : data_rom <= {16'd32605, 16'd3261};
                15'd15345 : data_rom <= {16'd32605, 16'd3258};
                15'd15346 : data_rom <= {16'd32605, 16'd3255};
                15'd15347 : data_rom <= {16'd32606, 16'd3252};
                15'd15348 : data_rom <= {16'd32606, 16'd3249};
                15'd15349 : data_rom <= {16'd32606, 16'd3246};
                15'd15350 : data_rom <= {16'd32607, 16'd3243};
                15'd15351 : data_rom <= {16'd32607, 16'd3240};
                15'd15352 : data_rom <= {16'd32607, 16'd3236};
                15'd15353 : data_rom <= {16'd32608, 16'd3233};
                15'd15354 : data_rom <= {16'd32608, 16'd3230};
                15'd15355 : data_rom <= {16'd32608, 16'd3227};
                15'd15356 : data_rom <= {16'd32608, 16'd3224};
                15'd15357 : data_rom <= {16'd32609, 16'd3221};
                15'd15358 : data_rom <= {16'd32609, 16'd3218};
                15'd15359 : data_rom <= {16'd32609, 16'd3214};
                15'd15360 : data_rom <= {16'd32610, 16'd3211};
                15'd15361 : data_rom <= {16'd32610, 16'd3208};
                15'd15362 : data_rom <= {16'd32610, 16'd3205};
                15'd15363 : data_rom <= {16'd32611, 16'd3202};
                15'd15364 : data_rom <= {16'd32611, 16'd3199};
                15'd15365 : data_rom <= {16'd32611, 16'd3196};
                15'd15366 : data_rom <= {16'd32612, 16'd3193};
                15'd15367 : data_rom <= {16'd32612, 16'd3189};
                15'd15368 : data_rom <= {16'd32612, 16'd3186};
                15'd15369 : data_rom <= {16'd32612, 16'd3183};
                15'd15370 : data_rom <= {16'd32613, 16'd3180};
                15'd15371 : data_rom <= {16'd32613, 16'd3177};
                15'd15372 : data_rom <= {16'd32613, 16'd3174};
                15'd15373 : data_rom <= {16'd32614, 16'd3171};
                15'd15374 : data_rom <= {16'd32614, 16'd3168};
                15'd15375 : data_rom <= {16'd32614, 16'd3164};
                15'd15376 : data_rom <= {16'd32615, 16'd3161};
                15'd15377 : data_rom <= {16'd32615, 16'd3158};
                15'd15378 : data_rom <= {16'd32615, 16'd3155};
                15'd15379 : data_rom <= {16'd32616, 16'd3152};
                15'd15380 : data_rom <= {16'd32616, 16'd3149};
                15'd15381 : data_rom <= {16'd32616, 16'd3146};
                15'd15382 : data_rom <= {16'd32616, 16'd3143};
                15'd15383 : data_rom <= {16'd32617, 16'd3139};
                15'd15384 : data_rom <= {16'd32617, 16'd3136};
                15'd15385 : data_rom <= {16'd32617, 16'd3133};
                15'd15386 : data_rom <= {16'd32618, 16'd3130};
                15'd15387 : data_rom <= {16'd32618, 16'd3127};
                15'd15388 : data_rom <= {16'd32618, 16'd3124};
                15'd15389 : data_rom <= {16'd32619, 16'd3121};
                15'd15390 : data_rom <= {16'd32619, 16'd3118};
                15'd15391 : data_rom <= {16'd32619, 16'd3114};
                15'd15392 : data_rom <= {16'd32619, 16'd3111};
                15'd15393 : data_rom <= {16'd32620, 16'd3108};
                15'd15394 : data_rom <= {16'd32620, 16'd3105};
                15'd15395 : data_rom <= {16'd32620, 16'd3102};
                15'd15396 : data_rom <= {16'd32621, 16'd3099};
                15'd15397 : data_rom <= {16'd32621, 16'd3096};
                15'd15398 : data_rom <= {16'd32621, 16'd3093};
                15'd15399 : data_rom <= {16'd32621, 16'd3089};
                15'd15400 : data_rom <= {16'd32622, 16'd3086};
                15'd15401 : data_rom <= {16'd32622, 16'd3083};
                15'd15402 : data_rom <= {16'd32622, 16'd3080};
                15'd15403 : data_rom <= {16'd32623, 16'd3077};
                15'd15404 : data_rom <= {16'd32623, 16'd3074};
                15'd15405 : data_rom <= {16'd32623, 16'd3071};
                15'd15406 : data_rom <= {16'd32624, 16'd3068};
                15'd15407 : data_rom <= {16'd32624, 16'd3064};
                15'd15408 : data_rom <= {16'd32624, 16'd3061};
                15'd15409 : data_rom <= {16'd32624, 16'd3058};
                15'd15410 : data_rom <= {16'd32625, 16'd3055};
                15'd15411 : data_rom <= {16'd32625, 16'd3052};
                15'd15412 : data_rom <= {16'd32625, 16'd3049};
                15'd15413 : data_rom <= {16'd32626, 16'd3046};
                15'd15414 : data_rom <= {16'd32626, 16'd3042};
                15'd15415 : data_rom <= {16'd32626, 16'd3039};
                15'd15416 : data_rom <= {16'd32626, 16'd3036};
                15'd15417 : data_rom <= {16'd32627, 16'd3033};
                15'd15418 : data_rom <= {16'd32627, 16'd3030};
                15'd15419 : data_rom <= {16'd32627, 16'd3027};
                15'd15420 : data_rom <= {16'd32628, 16'd3024};
                15'd15421 : data_rom <= {16'd32628, 16'd3021};
                15'd15422 : data_rom <= {16'd32628, 16'd3017};
                15'd15423 : data_rom <= {16'd32629, 16'd3014};
                15'd15424 : data_rom <= {16'd32629, 16'd3011};
                15'd15425 : data_rom <= {16'd32629, 16'd3008};
                15'd15426 : data_rom <= {16'd32629, 16'd3005};
                15'd15427 : data_rom <= {16'd32630, 16'd3002};
                15'd15428 : data_rom <= {16'd32630, 16'd2999};
                15'd15429 : data_rom <= {16'd32630, 16'd2996};
                15'd15430 : data_rom <= {16'd32631, 16'd2992};
                15'd15431 : data_rom <= {16'd32631, 16'd2989};
                15'd15432 : data_rom <= {16'd32631, 16'd2986};
                15'd15433 : data_rom <= {16'd32631, 16'd2983};
                15'd15434 : data_rom <= {16'd32632, 16'd2980};
                15'd15435 : data_rom <= {16'd32632, 16'd2977};
                15'd15436 : data_rom <= {16'd32632, 16'd2974};
                15'd15437 : data_rom <= {16'd32633, 16'd2971};
                15'd15438 : data_rom <= {16'd32633, 16'd2967};
                15'd15439 : data_rom <= {16'd32633, 16'd2964};
                15'd15440 : data_rom <= {16'd32633, 16'd2961};
                15'd15441 : data_rom <= {16'd32634, 16'd2958};
                15'd15442 : data_rom <= {16'd32634, 16'd2955};
                15'd15443 : data_rom <= {16'd32634, 16'd2952};
                15'd15444 : data_rom <= {16'd32635, 16'd2949};
                15'd15445 : data_rom <= {16'd32635, 16'd2946};
                15'd15446 : data_rom <= {16'd32635, 16'd2942};
                15'd15447 : data_rom <= {16'd32635, 16'd2939};
                15'd15448 : data_rom <= {16'd32636, 16'd2936};
                15'd15449 : data_rom <= {16'd32636, 16'd2933};
                15'd15450 : data_rom <= {16'd32636, 16'd2930};
                15'd15451 : data_rom <= {16'd32636, 16'd2927};
                15'd15452 : data_rom <= {16'd32637, 16'd2924};
                15'd15453 : data_rom <= {16'd32637, 16'd2920};
                15'd15454 : data_rom <= {16'd32637, 16'd2917};
                15'd15455 : data_rom <= {16'd32638, 16'd2914};
                15'd15456 : data_rom <= {16'd32638, 16'd2911};
                15'd15457 : data_rom <= {16'd32638, 16'd2908};
                15'd15458 : data_rom <= {16'd32638, 16'd2905};
                15'd15459 : data_rom <= {16'd32639, 16'd2902};
                15'd15460 : data_rom <= {16'd32639, 16'd2899};
                15'd15461 : data_rom <= {16'd32639, 16'd2895};
                15'd15462 : data_rom <= {16'd32640, 16'd2892};
                15'd15463 : data_rom <= {16'd32640, 16'd2889};
                15'd15464 : data_rom <= {16'd32640, 16'd2886};
                15'd15465 : data_rom <= {16'd32640, 16'd2883};
                15'd15466 : data_rom <= {16'd32641, 16'd2880};
                15'd15467 : data_rom <= {16'd32641, 16'd2877};
                15'd15468 : data_rom <= {16'd32641, 16'd2874};
                15'd15469 : data_rom <= {16'd32641, 16'd2870};
                15'd15470 : data_rom <= {16'd32642, 16'd2867};
                15'd15471 : data_rom <= {16'd32642, 16'd2864};
                15'd15472 : data_rom <= {16'd32642, 16'd2861};
                15'd15473 : data_rom <= {16'd32643, 16'd2858};
                15'd15474 : data_rom <= {16'd32643, 16'd2855};
                15'd15475 : data_rom <= {16'd32643, 16'd2852};
                15'd15476 : data_rom <= {16'd32643, 16'd2849};
                15'd15477 : data_rom <= {16'd32644, 16'd2845};
                15'd15478 : data_rom <= {16'd32644, 16'd2842};
                15'd15479 : data_rom <= {16'd32644, 16'd2839};
                15'd15480 : data_rom <= {16'd32645, 16'd2836};
                15'd15481 : data_rom <= {16'd32645, 16'd2833};
                15'd15482 : data_rom <= {16'd32645, 16'd2830};
                15'd15483 : data_rom <= {16'd32645, 16'd2827};
                15'd15484 : data_rom <= {16'd32646, 16'd2823};
                15'd15485 : data_rom <= {16'd32646, 16'd2820};
                15'd15486 : data_rom <= {16'd32646, 16'd2817};
                15'd15487 : data_rom <= {16'd32646, 16'd2814};
                15'd15488 : data_rom <= {16'd32647, 16'd2811};
                15'd15489 : data_rom <= {16'd32647, 16'd2808};
                15'd15490 : data_rom <= {16'd32647, 16'd2805};
                15'd15491 : data_rom <= {16'd32647, 16'd2802};
                15'd15492 : data_rom <= {16'd32648, 16'd2798};
                15'd15493 : data_rom <= {16'd32648, 16'd2795};
                15'd15494 : data_rom <= {16'd32648, 16'd2792};
                15'd15495 : data_rom <= {16'd32649, 16'd2789};
                15'd15496 : data_rom <= {16'd32649, 16'd2786};
                15'd15497 : data_rom <= {16'd32649, 16'd2783};
                15'd15498 : data_rom <= {16'd32649, 16'd2780};
                15'd15499 : data_rom <= {16'd32650, 16'd2777};
                15'd15500 : data_rom <= {16'd32650, 16'd2773};
                15'd15501 : data_rom <= {16'd32650, 16'd2770};
                15'd15502 : data_rom <= {16'd32650, 16'd2767};
                15'd15503 : data_rom <= {16'd32651, 16'd2764};
                15'd15504 : data_rom <= {16'd32651, 16'd2761};
                15'd15505 : data_rom <= {16'd32651, 16'd2758};
                15'd15506 : data_rom <= {16'd32651, 16'd2755};
                15'd15507 : data_rom <= {16'd32652, 16'd2751};
                15'd15508 : data_rom <= {16'd32652, 16'd2748};
                15'd15509 : data_rom <= {16'd32652, 16'd2745};
                15'd15510 : data_rom <= {16'd32653, 16'd2742};
                15'd15511 : data_rom <= {16'd32653, 16'd2739};
                15'd15512 : data_rom <= {16'd32653, 16'd2736};
                15'd15513 : data_rom <= {16'd32653, 16'd2733};
                15'd15514 : data_rom <= {16'd32654, 16'd2730};
                15'd15515 : data_rom <= {16'd32654, 16'd2726};
                15'd15516 : data_rom <= {16'd32654, 16'd2723};
                15'd15517 : data_rom <= {16'd32654, 16'd2720};
                15'd15518 : data_rom <= {16'd32655, 16'd2717};
                15'd15519 : data_rom <= {16'd32655, 16'd2714};
                15'd15520 : data_rom <= {16'd32655, 16'd2711};
                15'd15521 : data_rom <= {16'd32655, 16'd2708};
                15'd15522 : data_rom <= {16'd32656, 16'd2705};
                15'd15523 : data_rom <= {16'd32656, 16'd2701};
                15'd15524 : data_rom <= {16'd32656, 16'd2698};
                15'd15525 : data_rom <= {16'd32656, 16'd2695};
                15'd15526 : data_rom <= {16'd32657, 16'd2692};
                15'd15527 : data_rom <= {16'd32657, 16'd2689};
                15'd15528 : data_rom <= {16'd32657, 16'd2686};
                15'd15529 : data_rom <= {16'd32657, 16'd2683};
                15'd15530 : data_rom <= {16'd32658, 16'd2679};
                15'd15531 : data_rom <= {16'd32658, 16'd2676};
                15'd15532 : data_rom <= {16'd32658, 16'd2673};
                15'd15533 : data_rom <= {16'd32658, 16'd2670};
                15'd15534 : data_rom <= {16'd32659, 16'd2667};
                15'd15535 : data_rom <= {16'd32659, 16'd2664};
                15'd15536 : data_rom <= {16'd32659, 16'd2661};
                15'd15537 : data_rom <= {16'd32660, 16'd2658};
                15'd15538 : data_rom <= {16'd32660, 16'd2654};
                15'd15539 : data_rom <= {16'd32660, 16'd2651};
                15'd15540 : data_rom <= {16'd32660, 16'd2648};
                15'd15541 : data_rom <= {16'd32661, 16'd2645};
                15'd15542 : data_rom <= {16'd32661, 16'd2642};
                15'd15543 : data_rom <= {16'd32661, 16'd2639};
                15'd15544 : data_rom <= {16'd32661, 16'd2636};
                15'd15545 : data_rom <= {16'd32662, 16'd2633};
                15'd15546 : data_rom <= {16'd32662, 16'd2629};
                15'd15547 : data_rom <= {16'd32662, 16'd2626};
                15'd15548 : data_rom <= {16'd32662, 16'd2623};
                15'd15549 : data_rom <= {16'd32663, 16'd2620};
                15'd15550 : data_rom <= {16'd32663, 16'd2617};
                15'd15551 : data_rom <= {16'd32663, 16'd2614};
                15'd15552 : data_rom <= {16'd32663, 16'd2611};
                15'd15553 : data_rom <= {16'd32664, 16'd2607};
                15'd15554 : data_rom <= {16'd32664, 16'd2604};
                15'd15555 : data_rom <= {16'd32664, 16'd2601};
                15'd15556 : data_rom <= {16'd32664, 16'd2598};
                15'd15557 : data_rom <= {16'd32665, 16'd2595};
                15'd15558 : data_rom <= {16'd32665, 16'd2592};
                15'd15559 : data_rom <= {16'd32665, 16'd2589};
                15'd15560 : data_rom <= {16'd32665, 16'd2586};
                15'd15561 : data_rom <= {16'd32666, 16'd2582};
                15'd15562 : data_rom <= {16'd32666, 16'd2579};
                15'd15563 : data_rom <= {16'd32666, 16'd2576};
                15'd15564 : data_rom <= {16'd32666, 16'd2573};
                15'd15565 : data_rom <= {16'd32667, 16'd2570};
                15'd15566 : data_rom <= {16'd32667, 16'd2567};
                15'd15567 : data_rom <= {16'd32667, 16'd2564};
                15'd15568 : data_rom <= {16'd32667, 16'd2560};
                15'd15569 : data_rom <= {16'd32668, 16'd2557};
                15'd15570 : data_rom <= {16'd32668, 16'd2554};
                15'd15571 : data_rom <= {16'd32668, 16'd2551};
                15'd15572 : data_rom <= {16'd32668, 16'd2548};
                15'd15573 : data_rom <= {16'd32668, 16'd2545};
                15'd15574 : data_rom <= {16'd32669, 16'd2542};
                15'd15575 : data_rom <= {16'd32669, 16'd2539};
                15'd15576 : data_rom <= {16'd32669, 16'd2535};
                15'd15577 : data_rom <= {16'd32669, 16'd2532};
                15'd15578 : data_rom <= {16'd32670, 16'd2529};
                15'd15579 : data_rom <= {16'd32670, 16'd2526};
                15'd15580 : data_rom <= {16'd32670, 16'd2523};
                15'd15581 : data_rom <= {16'd32670, 16'd2520};
                15'd15582 : data_rom <= {16'd32671, 16'd2517};
                15'd15583 : data_rom <= {16'd32671, 16'd2513};
                15'd15584 : data_rom <= {16'd32671, 16'd2510};
                15'd15585 : data_rom <= {16'd32671, 16'd2507};
                15'd15586 : data_rom <= {16'd32672, 16'd2504};
                15'd15587 : data_rom <= {16'd32672, 16'd2501};
                15'd15588 : data_rom <= {16'd32672, 16'd2498};
                15'd15589 : data_rom <= {16'd32672, 16'd2495};
                15'd15590 : data_rom <= {16'd32673, 16'd2492};
                15'd15591 : data_rom <= {16'd32673, 16'd2488};
                15'd15592 : data_rom <= {16'd32673, 16'd2485};
                15'd15593 : data_rom <= {16'd32673, 16'd2482};
                15'd15594 : data_rom <= {16'd32674, 16'd2479};
                15'd15595 : data_rom <= {16'd32674, 16'd2476};
                15'd15596 : data_rom <= {16'd32674, 16'd2473};
                15'd15597 : data_rom <= {16'd32674, 16'd2470};
                15'd15598 : data_rom <= {16'd32675, 16'd2467};
                15'd15599 : data_rom <= {16'd32675, 16'd2463};
                15'd15600 : data_rom <= {16'd32675, 16'd2460};
                15'd15601 : data_rom <= {16'd32675, 16'd2457};
                15'd15602 : data_rom <= {16'd32675, 16'd2454};
                15'd15603 : data_rom <= {16'd32676, 16'd2451};
                15'd15604 : data_rom <= {16'd32676, 16'd2448};
                15'd15605 : data_rom <= {16'd32676, 16'd2445};
                15'd15606 : data_rom <= {16'd32676, 16'd2441};
                15'd15607 : data_rom <= {16'd32677, 16'd2438};
                15'd15608 : data_rom <= {16'd32677, 16'd2435};
                15'd15609 : data_rom <= {16'd32677, 16'd2432};
                15'd15610 : data_rom <= {16'd32677, 16'd2429};
                15'd15611 : data_rom <= {16'd32678, 16'd2426};
                15'd15612 : data_rom <= {16'd32678, 16'd2423};
                15'd15613 : data_rom <= {16'd32678, 16'd2420};
                15'd15614 : data_rom <= {16'd32678, 16'd2416};
                15'd15615 : data_rom <= {16'd32678, 16'd2413};
                15'd15616 : data_rom <= {16'd32679, 16'd2410};
                15'd15617 : data_rom <= {16'd32679, 16'd2407};
                15'd15618 : data_rom <= {16'd32679, 16'd2404};
                15'd15619 : data_rom <= {16'd32679, 16'd2401};
                15'd15620 : data_rom <= {16'd32680, 16'd2398};
                15'd15621 : data_rom <= {16'd32680, 16'd2394};
                15'd15622 : data_rom <= {16'd32680, 16'd2391};
                15'd15623 : data_rom <= {16'd32680, 16'd2388};
                15'd15624 : data_rom <= {16'd32681, 16'd2385};
                15'd15625 : data_rom <= {16'd32681, 16'd2382};
                15'd15626 : data_rom <= {16'd32681, 16'd2379};
                15'd15627 : data_rom <= {16'd32681, 16'd2376};
                15'd15628 : data_rom <= {16'd32681, 16'd2373};
                15'd15629 : data_rom <= {16'd32682, 16'd2369};
                15'd15630 : data_rom <= {16'd32682, 16'd2366};
                15'd15631 : data_rom <= {16'd32682, 16'd2363};
                15'd15632 : data_rom <= {16'd32682, 16'd2360};
                15'd15633 : data_rom <= {16'd32683, 16'd2357};
                15'd15634 : data_rom <= {16'd32683, 16'd2354};
                15'd15635 : data_rom <= {16'd32683, 16'd2351};
                15'd15636 : data_rom <= {16'd32683, 16'd2347};
                15'd15637 : data_rom <= {16'd32683, 16'd2344};
                15'd15638 : data_rom <= {16'd32684, 16'd2341};
                15'd15639 : data_rom <= {16'd32684, 16'd2338};
                15'd15640 : data_rom <= {16'd32684, 16'd2335};
                15'd15641 : data_rom <= {16'd32684, 16'd2332};
                15'd15642 : data_rom <= {16'd32685, 16'd2329};
                15'd15643 : data_rom <= {16'd32685, 16'd2326};
                15'd15644 : data_rom <= {16'd32685, 16'd2322};
                15'd15645 : data_rom <= {16'd32685, 16'd2319};
                15'd15646 : data_rom <= {16'd32686, 16'd2316};
                15'd15647 : data_rom <= {16'd32686, 16'd2313};
                15'd15648 : data_rom <= {16'd32686, 16'd2310};
                15'd15649 : data_rom <= {16'd32686, 16'd2307};
                15'd15650 : data_rom <= {16'd32686, 16'd2304};
                15'd15651 : data_rom <= {16'd32687, 16'd2300};
                15'd15652 : data_rom <= {16'd32687, 16'd2297};
                15'd15653 : data_rom <= {16'd32687, 16'd2294};
                15'd15654 : data_rom <= {16'd32687, 16'd2291};
                15'd15655 : data_rom <= {16'd32687, 16'd2288};
                15'd15656 : data_rom <= {16'd32688, 16'd2285};
                15'd15657 : data_rom <= {16'd32688, 16'd2282};
                15'd15658 : data_rom <= {16'd32688, 16'd2279};
                15'd15659 : data_rom <= {16'd32688, 16'd2275};
                15'd15660 : data_rom <= {16'd32689, 16'd2272};
                15'd15661 : data_rom <= {16'd32689, 16'd2269};
                15'd15662 : data_rom <= {16'd32689, 16'd2266};
                15'd15663 : data_rom <= {16'd32689, 16'd2263};
                15'd15664 : data_rom <= {16'd32689, 16'd2260};
                15'd15665 : data_rom <= {16'd32690, 16'd2257};
                15'd15666 : data_rom <= {16'd32690, 16'd2253};
                15'd15667 : data_rom <= {16'd32690, 16'd2250};
                15'd15668 : data_rom <= {16'd32690, 16'd2247};
                15'd15669 : data_rom <= {16'd32691, 16'd2244};
                15'd15670 : data_rom <= {16'd32691, 16'd2241};
                15'd15671 : data_rom <= {16'd32691, 16'd2238};
                15'd15672 : data_rom <= {16'd32691, 16'd2235};
                15'd15673 : data_rom <= {16'd32691, 16'd2231};
                15'd15674 : data_rom <= {16'd32692, 16'd2228};
                15'd15675 : data_rom <= {16'd32692, 16'd2225};
                15'd15676 : data_rom <= {16'd32692, 16'd2222};
                15'd15677 : data_rom <= {16'd32692, 16'd2219};
                15'd15678 : data_rom <= {16'd32692, 16'd2216};
                15'd15679 : data_rom <= {16'd32693, 16'd2213};
                15'd15680 : data_rom <= {16'd32693, 16'd2210};
                15'd15681 : data_rom <= {16'd32693, 16'd2206};
                15'd15682 : data_rom <= {16'd32693, 16'd2203};
                15'd15683 : data_rom <= {16'd32694, 16'd2200};
                15'd15684 : data_rom <= {16'd32694, 16'd2197};
                15'd15685 : data_rom <= {16'd32694, 16'd2194};
                15'd15686 : data_rom <= {16'd32694, 16'd2191};
                15'd15687 : data_rom <= {16'd32694, 16'd2188};
                15'd15688 : data_rom <= {16'd32695, 16'd2184};
                15'd15689 : data_rom <= {16'd32695, 16'd2181};
                15'd15690 : data_rom <= {16'd32695, 16'd2178};
                15'd15691 : data_rom <= {16'd32695, 16'd2175};
                15'd15692 : data_rom <= {16'd32695, 16'd2172};
                15'd15693 : data_rom <= {16'd32696, 16'd2169};
                15'd15694 : data_rom <= {16'd32696, 16'd2166};
                15'd15695 : data_rom <= {16'd32696, 16'd2163};
                15'd15696 : data_rom <= {16'd32696, 16'd2159};
                15'd15697 : data_rom <= {16'd32696, 16'd2156};
                15'd15698 : data_rom <= {16'd32697, 16'd2153};
                15'd15699 : data_rom <= {16'd32697, 16'd2150};
                15'd15700 : data_rom <= {16'd32697, 16'd2147};
                15'd15701 : data_rom <= {16'd32697, 16'd2144};
                15'd15702 : data_rom <= {16'd32697, 16'd2141};
                15'd15703 : data_rom <= {16'd32698, 16'd2137};
                15'd15704 : data_rom <= {16'd32698, 16'd2134};
                15'd15705 : data_rom <= {16'd32698, 16'd2131};
                15'd15706 : data_rom <= {16'd32698, 16'd2128};
                15'd15707 : data_rom <= {16'd32698, 16'd2125};
                15'd15708 : data_rom <= {16'd32699, 16'd2122};
                15'd15709 : data_rom <= {16'd32699, 16'd2119};
                15'd15710 : data_rom <= {16'd32699, 16'd2116};
                15'd15711 : data_rom <= {16'd32699, 16'd2112};
                15'd15712 : data_rom <= {16'd32700, 16'd2109};
                15'd15713 : data_rom <= {16'd32700, 16'd2106};
                15'd15714 : data_rom <= {16'd32700, 16'd2103};
                15'd15715 : data_rom <= {16'd32700, 16'd2100};
                15'd15716 : data_rom <= {16'd32700, 16'd2097};
                15'd15717 : data_rom <= {16'd32701, 16'd2094};
                15'd15718 : data_rom <= {16'd32701, 16'd2090};
                15'd15719 : data_rom <= {16'd32701, 16'd2087};
                15'd15720 : data_rom <= {16'd32701, 16'd2084};
                15'd15721 : data_rom <= {16'd32701, 16'd2081};
                15'd15722 : data_rom <= {16'd32702, 16'd2078};
                15'd15723 : data_rom <= {16'd32702, 16'd2075};
                15'd15724 : data_rom <= {16'd32702, 16'd2072};
                15'd15725 : data_rom <= {16'd32702, 16'd2068};
                15'd15726 : data_rom <= {16'd32702, 16'd2065};
                15'd15727 : data_rom <= {16'd32703, 16'd2062};
                15'd15728 : data_rom <= {16'd32703, 16'd2059};
                15'd15729 : data_rom <= {16'd32703, 16'd2056};
                15'd15730 : data_rom <= {16'd32703, 16'd2053};
                15'd15731 : data_rom <= {16'd32703, 16'd2050};
                15'd15732 : data_rom <= {16'd32703, 16'd2047};
                15'd15733 : data_rom <= {16'd32704, 16'd2043};
                15'd15734 : data_rom <= {16'd32704, 16'd2040};
                15'd15735 : data_rom <= {16'd32704, 16'd2037};
                15'd15736 : data_rom <= {16'd32704, 16'd2034};
                15'd15737 : data_rom <= {16'd32704, 16'd2031};
                15'd15738 : data_rom <= {16'd32705, 16'd2028};
                15'd15739 : data_rom <= {16'd32705, 16'd2025};
                15'd15740 : data_rom <= {16'd32705, 16'd2021};
                15'd15741 : data_rom <= {16'd32705, 16'd2018};
                15'd15742 : data_rom <= {16'd32705, 16'd2015};
                15'd15743 : data_rom <= {16'd32706, 16'd2012};
                15'd15744 : data_rom <= {16'd32706, 16'd2009};
                15'd15745 : data_rom <= {16'd32706, 16'd2006};
                15'd15746 : data_rom <= {16'd32706, 16'd2003};
                15'd15747 : data_rom <= {16'd32706, 16'd1999};
                15'd15748 : data_rom <= {16'd32707, 16'd1996};
                15'd15749 : data_rom <= {16'd32707, 16'd1993};
                15'd15750 : data_rom <= {16'd32707, 16'd1990};
                15'd15751 : data_rom <= {16'd32707, 16'd1987};
                15'd15752 : data_rom <= {16'd32707, 16'd1984};
                15'd15753 : data_rom <= {16'd32708, 16'd1981};
                15'd15754 : data_rom <= {16'd32708, 16'd1978};
                15'd15755 : data_rom <= {16'd32708, 16'd1974};
                15'd15756 : data_rom <= {16'd32708, 16'd1971};
                15'd15757 : data_rom <= {16'd32708, 16'd1968};
                15'd15758 : data_rom <= {16'd32708, 16'd1965};
                15'd15759 : data_rom <= {16'd32709, 16'd1962};
                15'd15760 : data_rom <= {16'd32709, 16'd1959};
                15'd15761 : data_rom <= {16'd32709, 16'd1956};
                15'd15762 : data_rom <= {16'd32709, 16'd1952};
                15'd15763 : data_rom <= {16'd32709, 16'd1949};
                15'd15764 : data_rom <= {16'd32710, 16'd1946};
                15'd15765 : data_rom <= {16'd32710, 16'd1943};
                15'd15766 : data_rom <= {16'd32710, 16'd1940};
                15'd15767 : data_rom <= {16'd32710, 16'd1937};
                15'd15768 : data_rom <= {16'd32710, 16'd1934};
                15'd15769 : data_rom <= {16'd32711, 16'd1931};
                15'd15770 : data_rom <= {16'd32711, 16'd1927};
                15'd15771 : data_rom <= {16'd32711, 16'd1924};
                15'd15772 : data_rom <= {16'd32711, 16'd1921};
                15'd15773 : data_rom <= {16'd32711, 16'd1918};
                15'd15774 : data_rom <= {16'd32711, 16'd1915};
                15'd15775 : data_rom <= {16'd32712, 16'd1912};
                15'd15776 : data_rom <= {16'd32712, 16'd1909};
                15'd15777 : data_rom <= {16'd32712, 16'd1905};
                15'd15778 : data_rom <= {16'd32712, 16'd1902};
                15'd15779 : data_rom <= {16'd32712, 16'd1899};
                15'd15780 : data_rom <= {16'd32713, 16'd1896};
                15'd15781 : data_rom <= {16'd32713, 16'd1893};
                15'd15782 : data_rom <= {16'd32713, 16'd1890};
                15'd15783 : data_rom <= {16'd32713, 16'd1887};
                15'd15784 : data_rom <= {16'd32713, 16'd1883};
                15'd15785 : data_rom <= {16'd32713, 16'd1880};
                15'd15786 : data_rom <= {16'd32714, 16'd1877};
                15'd15787 : data_rom <= {16'd32714, 16'd1874};
                15'd15788 : data_rom <= {16'd32714, 16'd1871};
                15'd15789 : data_rom <= {16'd32714, 16'd1868};
                15'd15790 : data_rom <= {16'd32714, 16'd1865};
                15'd15791 : data_rom <= {16'd32715, 16'd1862};
                15'd15792 : data_rom <= {16'd32715, 16'd1858};
                15'd15793 : data_rom <= {16'd32715, 16'd1855};
                15'd15794 : data_rom <= {16'd32715, 16'd1852};
                15'd15795 : data_rom <= {16'd32715, 16'd1849};
                15'd15796 : data_rom <= {16'd32715, 16'd1846};
                15'd15797 : data_rom <= {16'd32716, 16'd1843};
                15'd15798 : data_rom <= {16'd32716, 16'd1840};
                15'd15799 : data_rom <= {16'd32716, 16'd1836};
                15'd15800 : data_rom <= {16'd32716, 16'd1833};
                15'd15801 : data_rom <= {16'd32716, 16'd1830};
                15'd15802 : data_rom <= {16'd32716, 16'd1827};
                15'd15803 : data_rom <= {16'd32717, 16'd1824};
                15'd15804 : data_rom <= {16'd32717, 16'd1821};
                15'd15805 : data_rom <= {16'd32717, 16'd1818};
                15'd15806 : data_rom <= {16'd32717, 16'd1814};
                15'd15807 : data_rom <= {16'd32717, 16'd1811};
                15'd15808 : data_rom <= {16'd32718, 16'd1808};
                15'd15809 : data_rom <= {16'd32718, 16'd1805};
                15'd15810 : data_rom <= {16'd32718, 16'd1802};
                15'd15811 : data_rom <= {16'd32718, 16'd1799};
                15'd15812 : data_rom <= {16'd32718, 16'd1796};
                15'd15813 : data_rom <= {16'd32718, 16'd1793};
                15'd15814 : data_rom <= {16'd32719, 16'd1789};
                15'd15815 : data_rom <= {16'd32719, 16'd1786};
                15'd15816 : data_rom <= {16'd32719, 16'd1783};
                15'd15817 : data_rom <= {16'd32719, 16'd1780};
                15'd15818 : data_rom <= {16'd32719, 16'd1777};
                15'd15819 : data_rom <= {16'd32719, 16'd1774};
                15'd15820 : data_rom <= {16'd32720, 16'd1771};
                15'd15821 : data_rom <= {16'd32720, 16'd1767};
                15'd15822 : data_rom <= {16'd32720, 16'd1764};
                15'd15823 : data_rom <= {16'd32720, 16'd1761};
                15'd15824 : data_rom <= {16'd32720, 16'd1758};
                15'd15825 : data_rom <= {16'd32720, 16'd1755};
                15'd15826 : data_rom <= {16'd32721, 16'd1752};
                15'd15827 : data_rom <= {16'd32721, 16'd1749};
                15'd15828 : data_rom <= {16'd32721, 16'd1745};
                15'd15829 : data_rom <= {16'd32721, 16'd1742};
                15'd15830 : data_rom <= {16'd32721, 16'd1739};
                15'd15831 : data_rom <= {16'd32721, 16'd1736};
                15'd15832 : data_rom <= {16'd32722, 16'd1733};
                15'd15833 : data_rom <= {16'd32722, 16'd1730};
                15'd15834 : data_rom <= {16'd32722, 16'd1727};
                15'd15835 : data_rom <= {16'd32722, 16'd1723};
                15'd15836 : data_rom <= {16'd32722, 16'd1720};
                15'd15837 : data_rom <= {16'd32722, 16'd1717};
                15'd15838 : data_rom <= {16'd32723, 16'd1714};
                15'd15839 : data_rom <= {16'd32723, 16'd1711};
                15'd15840 : data_rom <= {16'd32723, 16'd1708};
                15'd15841 : data_rom <= {16'd32723, 16'd1705};
                15'd15842 : data_rom <= {16'd32723, 16'd1702};
                15'd15843 : data_rom <= {16'd32723, 16'd1698};
                15'd15844 : data_rom <= {16'd32724, 16'd1695};
                15'd15845 : data_rom <= {16'd32724, 16'd1692};
                15'd15846 : data_rom <= {16'd32724, 16'd1689};
                15'd15847 : data_rom <= {16'd32724, 16'd1686};
                15'd15848 : data_rom <= {16'd32724, 16'd1683};
                15'd15849 : data_rom <= {16'd32724, 16'd1680};
                15'd15850 : data_rom <= {16'd32725, 16'd1676};
                15'd15851 : data_rom <= {16'd32725, 16'd1673};
                15'd15852 : data_rom <= {16'd32725, 16'd1670};
                15'd15853 : data_rom <= {16'd32725, 16'd1667};
                15'd15854 : data_rom <= {16'd32725, 16'd1664};
                15'd15855 : data_rom <= {16'd32725, 16'd1661};
                15'd15856 : data_rom <= {16'd32726, 16'd1658};
                15'd15857 : data_rom <= {16'd32726, 16'd1654};
                15'd15858 : data_rom <= {16'd32726, 16'd1651};
                15'd15859 : data_rom <= {16'd32726, 16'd1648};
                15'd15860 : data_rom <= {16'd32726, 16'd1645};
                15'd15861 : data_rom <= {16'd32726, 16'd1642};
                15'd15862 : data_rom <= {16'd32726, 16'd1639};
                15'd15863 : data_rom <= {16'd32727, 16'd1636};
                15'd15864 : data_rom <= {16'd32727, 16'd1632};
                15'd15865 : data_rom <= {16'd32727, 16'd1629};
                15'd15866 : data_rom <= {16'd32727, 16'd1626};
                15'd15867 : data_rom <= {16'd32727, 16'd1623};
                15'd15868 : data_rom <= {16'd32727, 16'd1620};
                15'd15869 : data_rom <= {16'd32728, 16'd1617};
                15'd15870 : data_rom <= {16'd32728, 16'd1614};
                15'd15871 : data_rom <= {16'd32728, 16'd1611};
                15'd15872 : data_rom <= {16'd32728, 16'd1607};
                15'd15873 : data_rom <= {16'd32728, 16'd1604};
                15'd15874 : data_rom <= {16'd32728, 16'd1601};
                15'd15875 : data_rom <= {16'd32728, 16'd1598};
                15'd15876 : data_rom <= {16'd32729, 16'd1595};
                15'd15877 : data_rom <= {16'd32729, 16'd1592};
                15'd15878 : data_rom <= {16'd32729, 16'd1589};
                15'd15879 : data_rom <= {16'd32729, 16'd1585};
                15'd15880 : data_rom <= {16'd32729, 16'd1582};
                15'd15881 : data_rom <= {16'd32729, 16'd1579};
                15'd15882 : data_rom <= {16'd32730, 16'd1576};
                15'd15883 : data_rom <= {16'd32730, 16'd1573};
                15'd15884 : data_rom <= {16'd32730, 16'd1570};
                15'd15885 : data_rom <= {16'd32730, 16'd1567};
                15'd15886 : data_rom <= {16'd32730, 16'd1563};
                15'd15887 : data_rom <= {16'd32730, 16'd1560};
                15'd15888 : data_rom <= {16'd32730, 16'd1557};
                15'd15889 : data_rom <= {16'd32731, 16'd1554};
                15'd15890 : data_rom <= {16'd32731, 16'd1551};
                15'd15891 : data_rom <= {16'd32731, 16'd1548};
                15'd15892 : data_rom <= {16'd32731, 16'd1545};
                15'd15893 : data_rom <= {16'd32731, 16'd1541};
                15'd15894 : data_rom <= {16'd32731, 16'd1538};
                15'd15895 : data_rom <= {16'd32731, 16'd1535};
                15'd15896 : data_rom <= {16'd32732, 16'd1532};
                15'd15897 : data_rom <= {16'd32732, 16'd1529};
                15'd15898 : data_rom <= {16'd32732, 16'd1526};
                15'd15899 : data_rom <= {16'd32732, 16'd1523};
                15'd15900 : data_rom <= {16'd32732, 16'd1520};
                15'd15901 : data_rom <= {16'd32732, 16'd1516};
                15'd15902 : data_rom <= {16'd32733, 16'd1513};
                15'd15903 : data_rom <= {16'd32733, 16'd1510};
                15'd15904 : data_rom <= {16'd32733, 16'd1507};
                15'd15905 : data_rom <= {16'd32733, 16'd1504};
                15'd15906 : data_rom <= {16'd32733, 16'd1501};
                15'd15907 : data_rom <= {16'd32733, 16'd1498};
                15'd15908 : data_rom <= {16'd32733, 16'd1494};
                15'd15909 : data_rom <= {16'd32734, 16'd1491};
                15'd15910 : data_rom <= {16'd32734, 16'd1488};
                15'd15911 : data_rom <= {16'd32734, 16'd1485};
                15'd15912 : data_rom <= {16'd32734, 16'd1482};
                15'd15913 : data_rom <= {16'd32734, 16'd1479};
                15'd15914 : data_rom <= {16'd32734, 16'd1476};
                15'd15915 : data_rom <= {16'd32734, 16'd1472};
                15'd15916 : data_rom <= {16'd32735, 16'd1469};
                15'd15917 : data_rom <= {16'd32735, 16'd1466};
                15'd15918 : data_rom <= {16'd32735, 16'd1463};
                15'd15919 : data_rom <= {16'd32735, 16'd1460};
                15'd15920 : data_rom <= {16'd32735, 16'd1457};
                15'd15921 : data_rom <= {16'd32735, 16'd1454};
                15'd15922 : data_rom <= {16'd32735, 16'd1450};
                15'd15923 : data_rom <= {16'd32735, 16'd1447};
                15'd15924 : data_rom <= {16'd32736, 16'd1444};
                15'd15925 : data_rom <= {16'd32736, 16'd1441};
                15'd15926 : data_rom <= {16'd32736, 16'd1438};
                15'd15927 : data_rom <= {16'd32736, 16'd1435};
                15'd15928 : data_rom <= {16'd32736, 16'd1432};
                15'd15929 : data_rom <= {16'd32736, 16'd1429};
                15'd15930 : data_rom <= {16'd32736, 16'd1425};
                15'd15931 : data_rom <= {16'd32737, 16'd1422};
                15'd15932 : data_rom <= {16'd32737, 16'd1419};
                15'd15933 : data_rom <= {16'd32737, 16'd1416};
                15'd15934 : data_rom <= {16'd32737, 16'd1413};
                15'd15935 : data_rom <= {16'd32737, 16'd1410};
                15'd15936 : data_rom <= {16'd32737, 16'd1407};
                15'd15937 : data_rom <= {16'd32737, 16'd1403};
                15'd15938 : data_rom <= {16'd32738, 16'd1400};
                15'd15939 : data_rom <= {16'd32738, 16'd1397};
                15'd15940 : data_rom <= {16'd32738, 16'd1394};
                15'd15941 : data_rom <= {16'd32738, 16'd1391};
                15'd15942 : data_rom <= {16'd32738, 16'd1388};
                15'd15943 : data_rom <= {16'd32738, 16'd1385};
                15'd15944 : data_rom <= {16'd32738, 16'd1381};
                15'd15945 : data_rom <= {16'd32738, 16'd1378};
                15'd15946 : data_rom <= {16'd32739, 16'd1375};
                15'd15947 : data_rom <= {16'd32739, 16'd1372};
                15'd15948 : data_rom <= {16'd32739, 16'd1369};
                15'd15949 : data_rom <= {16'd32739, 16'd1366};
                15'd15950 : data_rom <= {16'd32739, 16'd1363};
                15'd15951 : data_rom <= {16'd32739, 16'd1359};
                15'd15952 : data_rom <= {16'd32739, 16'd1356};
                15'd15953 : data_rom <= {16'd32740, 16'd1353};
                15'd15954 : data_rom <= {16'd32740, 16'd1350};
                15'd15955 : data_rom <= {16'd32740, 16'd1347};
                15'd15956 : data_rom <= {16'd32740, 16'd1344};
                15'd15957 : data_rom <= {16'd32740, 16'd1341};
                15'd15958 : data_rom <= {16'd32740, 16'd1337};
                15'd15959 : data_rom <= {16'd32740, 16'd1334};
                15'd15960 : data_rom <= {16'd32740, 16'd1331};
                15'd15961 : data_rom <= {16'd32741, 16'd1328};
                15'd15962 : data_rom <= {16'd32741, 16'd1325};
                15'd15963 : data_rom <= {16'd32741, 16'd1322};
                15'd15964 : data_rom <= {16'd32741, 16'd1319};
                15'd15965 : data_rom <= {16'd32741, 16'd1316};
                15'd15966 : data_rom <= {16'd32741, 16'd1312};
                15'd15967 : data_rom <= {16'd32741, 16'd1309};
                15'd15968 : data_rom <= {16'd32741, 16'd1306};
                15'd15969 : data_rom <= {16'd32742, 16'd1303};
                15'd15970 : data_rom <= {16'd32742, 16'd1300};
                15'd15971 : data_rom <= {16'd32742, 16'd1297};
                15'd15972 : data_rom <= {16'd32742, 16'd1294};
                15'd15973 : data_rom <= {16'd32742, 16'd1290};
                15'd15974 : data_rom <= {16'd32742, 16'd1287};
                15'd15975 : data_rom <= {16'd32742, 16'd1284};
                15'd15976 : data_rom <= {16'd32742, 16'd1281};
                15'd15977 : data_rom <= {16'd32743, 16'd1278};
                15'd15978 : data_rom <= {16'd32743, 16'd1275};
                15'd15979 : data_rom <= {16'd32743, 16'd1272};
                15'd15980 : data_rom <= {16'd32743, 16'd1268};
                15'd15981 : data_rom <= {16'd32743, 16'd1265};
                15'd15982 : data_rom <= {16'd32743, 16'd1262};
                15'd15983 : data_rom <= {16'd32743, 16'd1259};
                15'd15984 : data_rom <= {16'd32743, 16'd1256};
                15'd15985 : data_rom <= {16'd32744, 16'd1253};
                15'd15986 : data_rom <= {16'd32744, 16'd1250};
                15'd15987 : data_rom <= {16'd32744, 16'd1246};
                15'd15988 : data_rom <= {16'd32744, 16'd1243};
                15'd15989 : data_rom <= {16'd32744, 16'd1240};
                15'd15990 : data_rom <= {16'd32744, 16'd1237};
                15'd15991 : data_rom <= {16'd32744, 16'd1234};
                15'd15992 : data_rom <= {16'd32744, 16'd1231};
                15'd15993 : data_rom <= {16'd32744, 16'd1228};
                15'd15994 : data_rom <= {16'd32745, 16'd1224};
                15'd15995 : data_rom <= {16'd32745, 16'd1221};
                15'd15996 : data_rom <= {16'd32745, 16'd1218};
                15'd15997 : data_rom <= {16'd32745, 16'd1215};
                15'd15998 : data_rom <= {16'd32745, 16'd1212};
                15'd15999 : data_rom <= {16'd32745, 16'd1209};
                15'd16000 : data_rom <= {16'd32745, 16'd1206};
                15'd16001 : data_rom <= {16'd32745, 16'd1203};
                15'd16002 : data_rom <= {16'd32746, 16'd1199};
                15'd16003 : data_rom <= {16'd32746, 16'd1196};
                15'd16004 : data_rom <= {16'd32746, 16'd1193};
                15'd16005 : data_rom <= {16'd32746, 16'd1190};
                15'd16006 : data_rom <= {16'd32746, 16'd1187};
                15'd16007 : data_rom <= {16'd32746, 16'd1184};
                15'd16008 : data_rom <= {16'd32746, 16'd1181};
                15'd16009 : data_rom <= {16'd32746, 16'd1177};
                15'd16010 : data_rom <= {16'd32746, 16'd1174};
                15'd16011 : data_rom <= {16'd32747, 16'd1171};
                15'd16012 : data_rom <= {16'd32747, 16'd1168};
                15'd16013 : data_rom <= {16'd32747, 16'd1165};
                15'd16014 : data_rom <= {16'd32747, 16'd1162};
                15'd16015 : data_rom <= {16'd32747, 16'd1159};
                15'd16016 : data_rom <= {16'd32747, 16'd1155};
                15'd16017 : data_rom <= {16'd32747, 16'd1152};
                15'd16018 : data_rom <= {16'd32747, 16'd1149};
                15'd16019 : data_rom <= {16'd32747, 16'd1146};
                15'd16020 : data_rom <= {16'd32748, 16'd1143};
                15'd16021 : data_rom <= {16'd32748, 16'd1140};
                15'd16022 : data_rom <= {16'd32748, 16'd1137};
                15'd16023 : data_rom <= {16'd32748, 16'd1133};
                15'd16024 : data_rom <= {16'd32748, 16'd1130};
                15'd16025 : data_rom <= {16'd32748, 16'd1127};
                15'd16026 : data_rom <= {16'd32748, 16'd1124};
                15'd16027 : data_rom <= {16'd32748, 16'd1121};
                15'd16028 : data_rom <= {16'd32748, 16'd1118};
                15'd16029 : data_rom <= {16'd32749, 16'd1115};
                15'd16030 : data_rom <= {16'd32749, 16'd1111};
                15'd16031 : data_rom <= {16'd32749, 16'd1108};
                15'd16032 : data_rom <= {16'd32749, 16'd1105};
                15'd16033 : data_rom <= {16'd32749, 16'd1102};
                15'd16034 : data_rom <= {16'd32749, 16'd1099};
                15'd16035 : data_rom <= {16'd32749, 16'd1096};
                15'd16036 : data_rom <= {16'd32749, 16'd1093};
                15'd16037 : data_rom <= {16'd32749, 16'd1089};
                15'd16038 : data_rom <= {16'd32749, 16'd1086};
                15'd16039 : data_rom <= {16'd32750, 16'd1083};
                15'd16040 : data_rom <= {16'd32750, 16'd1080};
                15'd16041 : data_rom <= {16'd32750, 16'd1077};
                15'd16042 : data_rom <= {16'd32750, 16'd1074};
                15'd16043 : data_rom <= {16'd32750, 16'd1071};
                15'd16044 : data_rom <= {16'd32750, 16'd1068};
                15'd16045 : data_rom <= {16'd32750, 16'd1064};
                15'd16046 : data_rom <= {16'd32750, 16'd1061};
                15'd16047 : data_rom <= {16'd32750, 16'd1058};
                15'd16048 : data_rom <= {16'd32750, 16'd1055};
                15'd16049 : data_rom <= {16'd32751, 16'd1052};
                15'd16050 : data_rom <= {16'd32751, 16'd1049};
                15'd16051 : data_rom <= {16'd32751, 16'd1046};
                15'd16052 : data_rom <= {16'd32751, 16'd1042};
                15'd16053 : data_rom <= {16'd32751, 16'd1039};
                15'd16054 : data_rom <= {16'd32751, 16'd1036};
                15'd16055 : data_rom <= {16'd32751, 16'd1033};
                15'd16056 : data_rom <= {16'd32751, 16'd1030};
                15'd16057 : data_rom <= {16'd32751, 16'd1027};
                15'd16058 : data_rom <= {16'd32751, 16'd1024};
                15'd16059 : data_rom <= {16'd32752, 16'd1020};
                15'd16060 : data_rom <= {16'd32752, 16'd1017};
                15'd16061 : data_rom <= {16'd32752, 16'd1014};
                15'd16062 : data_rom <= {16'd32752, 16'd1011};
                15'd16063 : data_rom <= {16'd32752, 16'd1008};
                15'd16064 : data_rom <= {16'd32752, 16'd1005};
                15'd16065 : data_rom <= {16'd32752, 16'd1002};
                15'd16066 : data_rom <= {16'd32752, 16'd998};
                15'd16067 : data_rom <= {16'd32752, 16'd995};
                15'd16068 : data_rom <= {16'd32752, 16'd992};
                15'd16069 : data_rom <= {16'd32753, 16'd989};
                15'd16070 : data_rom <= {16'd32753, 16'd986};
                15'd16071 : data_rom <= {16'd32753, 16'd983};
                15'd16072 : data_rom <= {16'd32753, 16'd980};
                15'd16073 : data_rom <= {16'd32753, 16'd976};
                15'd16074 : data_rom <= {16'd32753, 16'd973};
                15'd16075 : data_rom <= {16'd32753, 16'd970};
                15'd16076 : data_rom <= {16'd32753, 16'd967};
                15'd16077 : data_rom <= {16'd32753, 16'd964};
                15'd16078 : data_rom <= {16'd32753, 16'd961};
                15'd16079 : data_rom <= {16'd32753, 16'd958};
                15'd16080 : data_rom <= {16'd32754, 16'd954};
                15'd16081 : data_rom <= {16'd32754, 16'd951};
                15'd16082 : data_rom <= {16'd32754, 16'd948};
                15'd16083 : data_rom <= {16'd32754, 16'd945};
                15'd16084 : data_rom <= {16'd32754, 16'd942};
                15'd16085 : data_rom <= {16'd32754, 16'd939};
                15'd16086 : data_rom <= {16'd32754, 16'd936};
                15'd16087 : data_rom <= {16'd32754, 16'd932};
                15'd16088 : data_rom <= {16'd32754, 16'd929};
                15'd16089 : data_rom <= {16'd32754, 16'd926};
                15'd16090 : data_rom <= {16'd32754, 16'd923};
                15'd16091 : data_rom <= {16'd32755, 16'd920};
                15'd16092 : data_rom <= {16'd32755, 16'd917};
                15'd16093 : data_rom <= {16'd32755, 16'd914};
                15'd16094 : data_rom <= {16'd32755, 16'd910};
                15'd16095 : data_rom <= {16'd32755, 16'd907};
                15'd16096 : data_rom <= {16'd32755, 16'd904};
                15'd16097 : data_rom <= {16'd32755, 16'd901};
                15'd16098 : data_rom <= {16'd32755, 16'd898};
                15'd16099 : data_rom <= {16'd32755, 16'd895};
                15'd16100 : data_rom <= {16'd32755, 16'd892};
                15'd16101 : data_rom <= {16'd32755, 16'd889};
                15'd16102 : data_rom <= {16'd32756, 16'd885};
                15'd16103 : data_rom <= {16'd32756, 16'd882};
                15'd16104 : data_rom <= {16'd32756, 16'd879};
                15'd16105 : data_rom <= {16'd32756, 16'd876};
                15'd16106 : data_rom <= {16'd32756, 16'd873};
                15'd16107 : data_rom <= {16'd32756, 16'd870};
                15'd16108 : data_rom <= {16'd32756, 16'd867};
                15'd16109 : data_rom <= {16'd32756, 16'd863};
                15'd16110 : data_rom <= {16'd32756, 16'd860};
                15'd16111 : data_rom <= {16'd32756, 16'd857};
                15'd16112 : data_rom <= {16'd32756, 16'd854};
                15'd16113 : data_rom <= {16'd32756, 16'd851};
                15'd16114 : data_rom <= {16'd32757, 16'd848};
                15'd16115 : data_rom <= {16'd32757, 16'd845};
                15'd16116 : data_rom <= {16'd32757, 16'd841};
                15'd16117 : data_rom <= {16'd32757, 16'd838};
                15'd16118 : data_rom <= {16'd32757, 16'd835};
                15'd16119 : data_rom <= {16'd32757, 16'd832};
                15'd16120 : data_rom <= {16'd32757, 16'd829};
                15'd16121 : data_rom <= {16'd32757, 16'd826};
                15'd16122 : data_rom <= {16'd32757, 16'd823};
                15'd16123 : data_rom <= {16'd32757, 16'd819};
                15'd16124 : data_rom <= {16'd32757, 16'd816};
                15'd16125 : data_rom <= {16'd32757, 16'd813};
                15'd16126 : data_rom <= {16'd32757, 16'd810};
                15'd16127 : data_rom <= {16'd32758, 16'd807};
                15'd16128 : data_rom <= {16'd32758, 16'd804};
                15'd16129 : data_rom <= {16'd32758, 16'd801};
                15'd16130 : data_rom <= {16'd32758, 16'd797};
                15'd16131 : data_rom <= {16'd32758, 16'd794};
                15'd16132 : data_rom <= {16'd32758, 16'd791};
                15'd16133 : data_rom <= {16'd32758, 16'd788};
                15'd16134 : data_rom <= {16'd32758, 16'd785};
                15'd16135 : data_rom <= {16'd32758, 16'd782};
                15'd16136 : data_rom <= {16'd32758, 16'd779};
                15'd16137 : data_rom <= {16'd32758, 16'd775};
                15'd16138 : data_rom <= {16'd32758, 16'd772};
                15'd16139 : data_rom <= {16'd32758, 16'd769};
                15'd16140 : data_rom <= {16'd32759, 16'd766};
                15'd16141 : data_rom <= {16'd32759, 16'd763};
                15'd16142 : data_rom <= {16'd32759, 16'd760};
                15'd16143 : data_rom <= {16'd32759, 16'd757};
                15'd16144 : data_rom <= {16'd32759, 16'd753};
                15'd16145 : data_rom <= {16'd32759, 16'd750};
                15'd16146 : data_rom <= {16'd32759, 16'd747};
                15'd16147 : data_rom <= {16'd32759, 16'd744};
                15'd16148 : data_rom <= {16'd32759, 16'd741};
                15'd16149 : data_rom <= {16'd32759, 16'd738};
                15'd16150 : data_rom <= {16'd32759, 16'd735};
                15'd16151 : data_rom <= {16'd32759, 16'd731};
                15'd16152 : data_rom <= {16'd32759, 16'd728};
                15'd16153 : data_rom <= {16'd32759, 16'd725};
                15'd16154 : data_rom <= {16'd32760, 16'd722};
                15'd16155 : data_rom <= {16'd32760, 16'd719};
                15'd16156 : data_rom <= {16'd32760, 16'd716};
                15'd16157 : data_rom <= {16'd32760, 16'd713};
                15'd16158 : data_rom <= {16'd32760, 16'd709};
                15'd16159 : data_rom <= {16'd32760, 16'd706};
                15'd16160 : data_rom <= {16'd32760, 16'd703};
                15'd16161 : data_rom <= {16'd32760, 16'd700};
                15'd16162 : data_rom <= {16'd32760, 16'd697};
                15'd16163 : data_rom <= {16'd32760, 16'd694};
                15'd16164 : data_rom <= {16'd32760, 16'd691};
                15'd16165 : data_rom <= {16'd32760, 16'd688};
                15'd16166 : data_rom <= {16'd32760, 16'd684};
                15'd16167 : data_rom <= {16'd32760, 16'd681};
                15'd16168 : data_rom <= {16'd32760, 16'd678};
                15'd16169 : data_rom <= {16'd32761, 16'd675};
                15'd16170 : data_rom <= {16'd32761, 16'd672};
                15'd16171 : data_rom <= {16'd32761, 16'd669};
                15'd16172 : data_rom <= {16'd32761, 16'd666};
                15'd16173 : data_rom <= {16'd32761, 16'd662};
                15'd16174 : data_rom <= {16'd32761, 16'd659};
                15'd16175 : data_rom <= {16'd32761, 16'd656};
                15'd16176 : data_rom <= {16'd32761, 16'd653};
                15'd16177 : data_rom <= {16'd32761, 16'd650};
                15'd16178 : data_rom <= {16'd32761, 16'd647};
                15'd16179 : data_rom <= {16'd32761, 16'd644};
                15'd16180 : data_rom <= {16'd32761, 16'd640};
                15'd16181 : data_rom <= {16'd32761, 16'd637};
                15'd16182 : data_rom <= {16'd32761, 16'd634};
                15'd16183 : data_rom <= {16'd32761, 16'd631};
                15'd16184 : data_rom <= {16'd32761, 16'd628};
                15'd16185 : data_rom <= {16'd32762, 16'd625};
                15'd16186 : data_rom <= {16'd32762, 16'd622};
                15'd16187 : data_rom <= {16'd32762, 16'd618};
                15'd16188 : data_rom <= {16'd32762, 16'd615};
                15'd16189 : data_rom <= {16'd32762, 16'd612};
                15'd16190 : data_rom <= {16'd32762, 16'd609};
                15'd16191 : data_rom <= {16'd32762, 16'd606};
                15'd16192 : data_rom <= {16'd32762, 16'd603};
                15'd16193 : data_rom <= {16'd32762, 16'd600};
                15'd16194 : data_rom <= {16'd32762, 16'd596};
                15'd16195 : data_rom <= {16'd32762, 16'd593};
                15'd16196 : data_rom <= {16'd32762, 16'd590};
                15'd16197 : data_rom <= {16'd32762, 16'd587};
                15'd16198 : data_rom <= {16'd32762, 16'd584};
                15'd16199 : data_rom <= {16'd32762, 16'd581};
                15'd16200 : data_rom <= {16'd32762, 16'd578};
                15'd16201 : data_rom <= {16'd32762, 16'd574};
                15'd16202 : data_rom <= {16'd32763, 16'd571};
                15'd16203 : data_rom <= {16'd32763, 16'd568};
                15'd16204 : data_rom <= {16'd32763, 16'd565};
                15'd16205 : data_rom <= {16'd32763, 16'd562};
                15'd16206 : data_rom <= {16'd32763, 16'd559};
                15'd16207 : data_rom <= {16'd32763, 16'd556};
                15'd16208 : data_rom <= {16'd32763, 16'd552};
                15'd16209 : data_rom <= {16'd32763, 16'd549};
                15'd16210 : data_rom <= {16'd32763, 16'd546};
                15'd16211 : data_rom <= {16'd32763, 16'd543};
                15'd16212 : data_rom <= {16'd32763, 16'd540};
                15'd16213 : data_rom <= {16'd32763, 16'd537};
                15'd16214 : data_rom <= {16'd32763, 16'd534};
                15'd16215 : data_rom <= {16'd32763, 16'd530};
                15'd16216 : data_rom <= {16'd32763, 16'd527};
                15'd16217 : data_rom <= {16'd32763, 16'd524};
                15'd16218 : data_rom <= {16'd32763, 16'd521};
                15'd16219 : data_rom <= {16'd32763, 16'd518};
                15'd16220 : data_rom <= {16'd32763, 16'd515};
                15'd16221 : data_rom <= {16'd32763, 16'd512};
                15'd16222 : data_rom <= {16'd32764, 16'd508};
                15'd16223 : data_rom <= {16'd32764, 16'd505};
                15'd16224 : data_rom <= {16'd32764, 16'd502};
                15'd16225 : data_rom <= {16'd32764, 16'd499};
                15'd16226 : data_rom <= {16'd32764, 16'd496};
                15'd16227 : data_rom <= {16'd32764, 16'd493};
                15'd16228 : data_rom <= {16'd32764, 16'd490};
                15'd16229 : data_rom <= {16'd32764, 16'd486};
                15'd16230 : data_rom <= {16'd32764, 16'd483};
                15'd16231 : data_rom <= {16'd32764, 16'd480};
                15'd16232 : data_rom <= {16'd32764, 16'd477};
                15'd16233 : data_rom <= {16'd32764, 16'd474};
                15'd16234 : data_rom <= {16'd32764, 16'd471};
                15'd16235 : data_rom <= {16'd32764, 16'd468};
                15'd16236 : data_rom <= {16'd32764, 16'd464};
                15'd16237 : data_rom <= {16'd32764, 16'd461};
                15'd16238 : data_rom <= {16'd32764, 16'd458};
                15'd16239 : data_rom <= {16'd32764, 16'd455};
                15'd16240 : data_rom <= {16'd32764, 16'd452};
                15'd16241 : data_rom <= {16'd32764, 16'd449};
                15'd16242 : data_rom <= {16'd32764, 16'd446};
                15'd16243 : data_rom <= {16'd32765, 16'd442};
                15'd16244 : data_rom <= {16'd32765, 16'd439};
                15'd16245 : data_rom <= {16'd32765, 16'd436};
                15'd16246 : data_rom <= {16'd32765, 16'd433};
                15'd16247 : data_rom <= {16'd32765, 16'd430};
                15'd16248 : data_rom <= {16'd32765, 16'd427};
                15'd16249 : data_rom <= {16'd32765, 16'd424};
                15'd16250 : data_rom <= {16'd32765, 16'd421};
                15'd16251 : data_rom <= {16'd32765, 16'd417};
                15'd16252 : data_rom <= {16'd32765, 16'd414};
                15'd16253 : data_rom <= {16'd32765, 16'd411};
                15'd16254 : data_rom <= {16'd32765, 16'd408};
                15'd16255 : data_rom <= {16'd32765, 16'd405};
                15'd16256 : data_rom <= {16'd32765, 16'd402};
                15'd16257 : data_rom <= {16'd32765, 16'd399};
                15'd16258 : data_rom <= {16'd32765, 16'd395};
                15'd16259 : data_rom <= {16'd32765, 16'd392};
                15'd16260 : data_rom <= {16'd32765, 16'd389};
                15'd16261 : data_rom <= {16'd32765, 16'd386};
                15'd16262 : data_rom <= {16'd32765, 16'd383};
                15'd16263 : data_rom <= {16'd32765, 16'd380};
                15'd16264 : data_rom <= {16'd32765, 16'd377};
                15'd16265 : data_rom <= {16'd32765, 16'd373};
                15'd16266 : data_rom <= {16'd32765, 16'd370};
                15'd16267 : data_rom <= {16'd32765, 16'd367};
                15'd16268 : data_rom <= {16'd32765, 16'd364};
                15'd16269 : data_rom <= {16'd32766, 16'd361};
                15'd16270 : data_rom <= {16'd32766, 16'd358};
                15'd16271 : data_rom <= {16'd32766, 16'd355};
                15'd16272 : data_rom <= {16'd32766, 16'd351};
                15'd16273 : data_rom <= {16'd32766, 16'd348};
                15'd16274 : data_rom <= {16'd32766, 16'd345};
                15'd16275 : data_rom <= {16'd32766, 16'd342};
                15'd16276 : data_rom <= {16'd32766, 16'd339};
                15'd16277 : data_rom <= {16'd32766, 16'd336};
                15'd16278 : data_rom <= {16'd32766, 16'd333};
                15'd16279 : data_rom <= {16'd32766, 16'd329};
                15'd16280 : data_rom <= {16'd32766, 16'd326};
                15'd16281 : data_rom <= {16'd32766, 16'd323};
                15'd16282 : data_rom <= {16'd32766, 16'd320};
                15'd16283 : data_rom <= {16'd32766, 16'd317};
                15'd16284 : data_rom <= {16'd32766, 16'd314};
                15'd16285 : data_rom <= {16'd32766, 16'd311};
                15'd16286 : data_rom <= {16'd32766, 16'd307};
                15'd16287 : data_rom <= {16'd32766, 16'd304};
                15'd16288 : data_rom <= {16'd32766, 16'd301};
                15'd16289 : data_rom <= {16'd32766, 16'd298};
                15'd16290 : data_rom <= {16'd32766, 16'd295};
                15'd16291 : data_rom <= {16'd32766, 16'd292};
                15'd16292 : data_rom <= {16'd32766, 16'd289};
                15'd16293 : data_rom <= {16'd32766, 16'd285};
                15'd16294 : data_rom <= {16'd32766, 16'd282};
                15'd16295 : data_rom <= {16'd32766, 16'd279};
                15'd16296 : data_rom <= {16'd32766, 16'd276};
                15'd16297 : data_rom <= {16'd32766, 16'd273};
                15'd16298 : data_rom <= {16'd32766, 16'd270};
                15'd16299 : data_rom <= {16'd32766, 16'd267};
                15'd16300 : data_rom <= {16'd32766, 16'd263};
                15'd16301 : data_rom <= {16'd32766, 16'd260};
                15'd16302 : data_rom <= {16'd32766, 16'd257};
                15'd16303 : data_rom <= {16'd32767, 16'd254};
                15'd16304 : data_rom <= {16'd32767, 16'd251};
                15'd16305 : data_rom <= {16'd32767, 16'd248};
                15'd16306 : data_rom <= {16'd32767, 16'd245};
                15'd16307 : data_rom <= {16'd32767, 16'd241};
                15'd16308 : data_rom <= {16'd32767, 16'd238};
                15'd16309 : data_rom <= {16'd32767, 16'd235};
                15'd16310 : data_rom <= {16'd32767, 16'd232};
                15'd16311 : data_rom <= {16'd32767, 16'd229};
                15'd16312 : data_rom <= {16'd32767, 16'd226};
                15'd16313 : data_rom <= {16'd32767, 16'd223};
                15'd16314 : data_rom <= {16'd32767, 16'd219};
                15'd16315 : data_rom <= {16'd32767, 16'd216};
                15'd16316 : data_rom <= {16'd32767, 16'd213};
                15'd16317 : data_rom <= {16'd32767, 16'd210};
                15'd16318 : data_rom <= {16'd32767, 16'd207};
                15'd16319 : data_rom <= {16'd32767, 16'd204};
                15'd16320 : data_rom <= {16'd32767, 16'd201};
                15'd16321 : data_rom <= {16'd32767, 16'd197};
                15'd16322 : data_rom <= {16'd32767, 16'd194};
                15'd16323 : data_rom <= {16'd32767, 16'd191};
                15'd16324 : data_rom <= {16'd32767, 16'd188};
                15'd16325 : data_rom <= {16'd32767, 16'd185};
                15'd16326 : data_rom <= {16'd32767, 16'd182};
                15'd16327 : data_rom <= {16'd32767, 16'd179};
                15'd16328 : data_rom <= {16'd32767, 16'd175};
                15'd16329 : data_rom <= {16'd32767, 16'd172};
                15'd16330 : data_rom <= {16'd32767, 16'd169};
                15'd16331 : data_rom <= {16'd32767, 16'd166};
                15'd16332 : data_rom <= {16'd32767, 16'd163};
                15'd16333 : data_rom <= {16'd32767, 16'd160};
                15'd16334 : data_rom <= {16'd32767, 16'd157};
                15'd16335 : data_rom <= {16'd32767, 16'd153};
                15'd16336 : data_rom <= {16'd32767, 16'd150};
                15'd16337 : data_rom <= {16'd32767, 16'd147};
                15'd16338 : data_rom <= {16'd32767, 16'd144};
                15'd16339 : data_rom <= {16'd32767, 16'd141};
                15'd16340 : data_rom <= {16'd32767, 16'd138};
                15'd16341 : data_rom <= {16'd32767, 16'd135};
                15'd16342 : data_rom <= {16'd32767, 16'd131};
                15'd16343 : data_rom <= {16'd32767, 16'd128};
                15'd16344 : data_rom <= {16'd32767, 16'd125};
                15'd16345 : data_rom <= {16'd32767, 16'd122};
                15'd16346 : data_rom <= {16'd32767, 16'd119};
                15'd16347 : data_rom <= {16'd32767, 16'd116};
                15'd16348 : data_rom <= {16'd32767, 16'd113};
                15'd16349 : data_rom <= {16'd32767, 16'd110};
                15'd16350 : data_rom <= {16'd32767, 16'd106};
                15'd16351 : data_rom <= {16'd32767, 16'd103};
                15'd16352 : data_rom <= {16'd32767, 16'd100};
                15'd16353 : data_rom <= {16'd32767, 16'd97};
                15'd16354 : data_rom <= {16'd32767, 16'd94};
                15'd16355 : data_rom <= {16'd32767, 16'd91};
                15'd16356 : data_rom <= {16'd32767, 16'd88};
                15'd16357 : data_rom <= {16'd32767, 16'd84};
                15'd16358 : data_rom <= {16'd32767, 16'd81};
                15'd16359 : data_rom <= {16'd32767, 16'd78};
                15'd16360 : data_rom <= {16'd32767, 16'd75};
                15'd16361 : data_rom <= {16'd32767, 16'd72};
                15'd16362 : data_rom <= {16'd32767, 16'd69};
                15'd16363 : data_rom <= {16'd32767, 16'd66};
                15'd16364 : data_rom <= {16'd32767, 16'd62};
                15'd16365 : data_rom <= {16'd32767, 16'd59};
                15'd16366 : data_rom <= {16'd32767, 16'd56};
                15'd16367 : data_rom <= {16'd32767, 16'd53};
                15'd16368 : data_rom <= {16'd32767, 16'd50};
                15'd16369 : data_rom <= {16'd32767, 16'd47};
                15'd16370 : data_rom <= {16'd32767, 16'd44};
                15'd16371 : data_rom <= {16'd32767, 16'd40};
                15'd16372 : data_rom <= {16'd32767, 16'd37};
                15'd16373 : data_rom <= {16'd32767, 16'd34};
                15'd16374 : data_rom <= {16'd32767, 16'd31};
                15'd16375 : data_rom <= {16'd32767, 16'd28};
                15'd16376 : data_rom <= {16'd32767, 16'd25};
                15'd16377 : data_rom <= {16'd32767, 16'd22};
                15'd16378 : data_rom <= {16'd32767, 16'd18};
                15'd16379 : data_rom <= {16'd32767, 16'd15};
                15'd16380 : data_rom <= {16'd32767, 16'd12};
                15'd16381 : data_rom <= {16'd32767, 16'd9};
                15'd16382 : data_rom <= {16'd32767, 16'd6};
                15'd16383 : data_rom <= {16'd32767, 16'd3};
				default : data_rom <= 32'hABCDEFAB;				
			endcase
		end
	
	//n사분면 bit에 따라 data_rom의 부호 조절
	always @ (*)
		begin
			case(addr[15:14])
				2'b00 : begin
					sin_out <= data_rom[31:16];
					cos_out <= data_rom[15:0];
					end
				2'b01 : begin
					sin_out <= data_rom[31:16];
					cos_out <= (~data_rom[15:0] + 2);
					end
				2'b10 : begin
					sin_out <= (~data_rom[31:16] +2);
					cos_out <= (~data_rom[15:0] + 2);
					end
				2'b11 : begin
					sin_out <= (~data_rom[31:16] +2);
					cos_out <= data_rom[15:0];
					end
				default : begin
					sin_out <= (~data_rom[31:16] +2);
					cos_out <= data_rom[15:0];
					end
			endcase
		end
endmodule
